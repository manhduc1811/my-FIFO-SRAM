/************************************************************************************************
************************************************************************************************/
module mySRAM_tb;
    parameter       BITS = 12, WORD_DEPTH = 1024, ADDR_WIDTH = 10;
    reg             clk,rst_n;
    reg             read;
    reg             write;
    reg  [BITS-1:0] data_in;
    wire [BITS-1:0] data_out;
    wire            ready;
    wire            overflow;
    mySRAM #(
		.BITS(BITS),
		.WORD_DEPTH(WORD_DEPTH),
		.ADDR_WIDTH(ADDR_WIDTH)
	) 
	UUT (
		.clk(clk),
		.rst_n(rst_n),
		.read(read),
		.write(write),
		.data_in(data_in),
		.data_out(data_out),
		.ready(ready),
		.overflow(overflow)
	);
    always #10 clk  = !clk;
    initial begin
            clk     = 0;
            rst_n   = 0;
            read    = 0;
            write   = 0;
        #20 rst_n   = 1;
			data_in = 12'h000;		write   = 1;		
        #20 data_in = 12'h001; 
        #20 data_in = 12'h002; 
        #20 data_in = 12'h003; 
        #20 data_in = 12'h004; 
        #20 data_in = 12'h005;		read    = 1;		
        #20 data_in = 12'h006; 
        #20 data_in = 12'h007; 
        #20 data_in = 12'h008; 		read    = 0;
        #20 data_in = 12'h009; 
        #20 data_in = 12'h00a; 
        #20 data_in = 12'h00b; 
        #20 data_in = 12'h00c; 
        #20 data_in = 12'h00d; 
        #20 data_in = 12'h00e; 
        #20 data_in = 12'h00f; 
        #20 data_in = 12'h010; 
        #20 data_in = 12'h011; 
        #20 data_in = 12'h012; 
        #20 data_in = 12'h013; 
        #20 data_in = 12'h014; 
        #20 data_in = 12'h015; 
        #20 data_in = 12'h016; 
        #20 data_in = 12'h017; 
        #20 data_in = 12'h018; 
        #20 data_in = 12'h019; 
        #20 data_in = 12'h01a; 
        #20 data_in = 12'h01b; 
        #20 data_in = 12'h01c; 
        #20 data_in = 12'h01d; 
        #20 data_in = 12'h01e; 
        #20 data_in = 12'h01f; 
        #20 data_in = 12'h020; 
        #20 data_in = 12'h021; 
        #20 data_in = 12'h022; 
        #20 data_in = 12'h023; 
        #20 data_in = 12'h024; 
        #20 data_in = 12'h025; 
        #20 data_in = 12'h026; 
        #20 data_in = 12'h027; 
        #20 data_in = 12'h028; 
        #20 data_in = 12'h029; 
        #20 data_in = 12'h02a; 
        #20 data_in = 12'h02b; 
        #20 data_in = 12'h02c; 
        #20 data_in = 12'h02d; 
        #20 data_in = 12'h02e; 
        #20 data_in = 12'h02f; 
        #20 data_in = 12'h030; 
        #20 data_in = 12'h031; 
        #20 data_in = 12'h032; 
        #20 data_in = 12'h033; 
        #20 data_in = 12'h034; 
        #20 data_in = 12'h035; 
        #20 data_in = 12'h036; 
        #20 data_in = 12'h037; 
        #20 data_in = 12'h038; 
        #20 data_in = 12'h039; 
        #20 data_in = 12'h03a; 
        #20 data_in = 12'h03b; 
        #20 data_in = 12'h03c; 
        #20 data_in = 12'h03d; 
        #20 data_in = 12'h03e; 
        #20 data_in = 12'h03f; 
        #20 data_in = 12'h040; 
        #20 data_in = 12'h041; 
        #20 data_in = 12'h042; 
        #20 data_in = 12'h043; 
        #20 data_in = 12'h044; 
        #20 data_in = 12'h045; 
        #20 data_in = 12'h046; 
        #20 data_in = 12'h047; 
        #20 data_in = 12'h048; 
        #20 data_in = 12'h049; 
        #20 data_in = 12'h04a; 
        #20 data_in = 12'h04b; 
        #20 data_in = 12'h04c; 
        #20 data_in = 12'h04d; 
        #20 data_in = 12'h04e; 
        #20 data_in = 12'h04f; 
        #20 data_in = 12'h050; 
        #20 data_in = 12'h051; 
        #20 data_in = 12'h052; 
        #20 data_in = 12'h053; 
        #20 data_in = 12'h054; 
        #20 data_in = 12'h055; 
        #20 data_in = 12'h056; 
        #20 data_in = 12'h057; 
        #20 data_in = 12'h058; 
        #20 data_in = 12'h059; 
        #20 data_in = 12'h05a; 
        #20 data_in = 12'h05b; 
        #20 data_in = 12'h05c; 
        #20 data_in = 12'h05d; 
        #20 data_in = 12'h05e; 
        #20 data_in = 12'h05f; 
        #20 data_in = 12'h060; 
        #20 data_in = 12'h061; 
        #20 data_in = 12'h062; 
        #20 data_in = 12'h063; 
        #20 data_in = 12'h064; 
        #20 data_in = 12'h065; 
        #20 data_in = 12'h066; 
        #20 data_in = 12'h067; 
        #20 data_in = 12'h068; 
        #20 data_in = 12'h069; 
        #20 data_in = 12'h06a; 
        #20 data_in = 12'h06b; 
        #20 data_in = 12'h06c; 
        #20 data_in = 12'h06d; 
        #20 data_in = 12'h06e; 
        #20 data_in = 12'h06f; 
        #20 data_in = 12'h070; 
        #20 data_in = 12'h071; 
        #20 data_in = 12'h072; 
        #20 data_in = 12'h073; 
        #20 data_in = 12'h074; 
        #20 data_in = 12'h075; 
        #20 data_in = 12'h076; 
        #20 data_in = 12'h077; 
        #20 data_in = 12'h078; 
        #20 data_in = 12'h079; 
        #20 data_in = 12'h07a; 
        #20 data_in = 12'h07b; 
        #20 data_in = 12'h07c; 
        #20 data_in = 12'h07d; 
        #20 data_in = 12'h07e; 
        #20 data_in = 12'h07f; 
        #20 data_in = 12'h080; 
        #20 data_in = 12'h081; 
        #20 data_in = 12'h082; 
        #20 data_in = 12'h083; 
        #20 data_in = 12'h084; 
        #20 data_in = 12'h085; 
        #20 data_in = 12'h086; 
        #20 data_in = 12'h087; 
        #20 data_in = 12'h088; 
        #20 data_in = 12'h089; 
        #20 data_in = 12'h08a; 
        #20 data_in = 12'h08b; 
        #20 data_in = 12'h08c; 
        #20 data_in = 12'h08d; 
        #20 data_in = 12'h08e; 
        #20 data_in = 12'h08f; 
        #20 data_in = 12'h090; 
        #20 data_in = 12'h091; 
        #20 data_in = 12'h092; 
        #20 data_in = 12'h093; 
        #20 data_in = 12'h094; 
        #20 data_in = 12'h095; 
        #20 data_in = 12'h096; 
        #20 data_in = 12'h097; 
        #20 data_in = 12'h098; 
        #20 data_in = 12'h099; 
        #20 data_in = 12'h09a; 
        #20 data_in = 12'h09b; 
        #20 data_in = 12'h09c; 
        #20 data_in = 12'h09d; 
        #20 data_in = 12'h09e; 
        #20 data_in = 12'h09f; 
        #20 data_in = 12'h0a0; 
        #20 data_in = 12'h0a1; 
        #20 data_in = 12'h0a2; 
        #20 data_in = 12'h0a3; 
        #20 data_in = 12'h0a4; 
        #20 data_in = 12'h0a5; 
        #20 data_in = 12'h0a6; 
        #20 data_in = 12'h0a7; 
        #20 data_in = 12'h0a8; 
        #20 data_in = 12'h0a9; 
        #20 data_in = 12'h0aa; 
        #20 data_in = 12'h0ab; 
        #20 data_in = 12'h0ac; 
        #20 data_in = 12'h0ad; 
        #20 data_in = 12'h0ae; 
        #20 data_in = 12'h0af; 
        #20 data_in = 12'h0b0; 
        #20 data_in = 12'h0b1; 
        #20 data_in = 12'h0b2; 
        #20 data_in = 12'h0b3; 
        #20 data_in = 12'h0b4; 
        #20 data_in = 12'h0b5; 
        #20 data_in = 12'h0b6; 
        #20 data_in = 12'h0b7; 
        #20 data_in = 12'h0b8; 
        #20 data_in = 12'h0b9; 
        #20 data_in = 12'h0ba; 
        #20 data_in = 12'h0bb; 
        #20 data_in = 12'h0bc; 
        #20 data_in = 12'h0bd; 
        #20 data_in = 12'h0be; 
        #20 data_in = 12'h0bf; 
        #20 data_in = 12'h0c0; 
        #20 data_in = 12'h0c1; 
        #20 data_in = 12'h0c2; 
        #20 data_in = 12'h0c3; 
        #20 data_in = 12'h0c4; 
        #20 data_in = 12'h0c5; 
        #20 data_in = 12'h0c6; 
        #20 data_in = 12'h0c7; 
        #20 data_in = 12'h0c8; 
        #20 data_in = 12'h0c9; 
        #20 data_in = 12'h0ca; 
        #20 data_in = 12'h0cb; 
        #20 data_in = 12'h0cc; 
        #20 data_in = 12'h0cd; 
        #20 data_in = 12'h0ce; 
        #20 data_in = 12'h0cf; 
        #20 data_in = 12'h0d0; 
        #20 data_in = 12'h0d1; 
        #20 data_in = 12'h0d2; 
        #20 data_in = 12'h0d3; 
        #20 data_in = 12'h0d4; 
        #20 data_in = 12'h0d5; 
        #20 data_in = 12'h0d6; 
        #20 data_in = 12'h0d7; 
        #20 data_in = 12'h0d8; 
        #20 data_in = 12'h0d9; 
        #20 data_in = 12'h0da; 
        #20 data_in = 12'h0db; 
        #20 data_in = 12'h0dc; 
        #20 data_in = 12'h0dd; 
        #20 data_in = 12'h0de; 
        #20 data_in = 12'h0df; 
        #20 data_in = 12'h0e0; 
        #20 data_in = 12'h0e1; 
        #20 data_in = 12'h0e2; 
        #20 data_in = 12'h0e3; 
        #20 data_in = 12'h0e4; 
        #20 data_in = 12'h0e5; 
        #20 data_in = 12'h0e6; 
        #20 data_in = 12'h0e7; 
        #20 data_in = 12'h0e8; 
        #20 data_in = 12'h0e9; 
        #20 data_in = 12'h0ea; 
        #20 data_in = 12'h0eb; 
        #20 data_in = 12'h0ec; 
        #20 data_in = 12'h0ed; 
        #20 data_in = 12'h0ee; 
        #20 data_in = 12'h0ef; 
        #20 data_in = 12'h0f0; 
        #20 data_in = 12'h0f1; 
        #20 data_in = 12'h0f2; 
        #20 data_in = 12'h0f3; 
        #20 data_in = 12'h0f4; 
        #20 data_in = 12'h0f5; 
        #20 data_in = 12'h0f6; 
        #20 data_in = 12'h0f7; 
        #20 data_in = 12'h0f8; 
        #20 data_in = 12'h0f9; 
        #20 data_in = 12'h0fa; 
        #20 data_in = 12'h0fb; 
        #20 data_in = 12'h0fc; 
        #20 data_in = 12'h0fd; 
        #20 data_in = 12'h0fe; 
        #20 data_in = 12'h0ff; 
        #20 data_in = 12'h100; 
        #20 data_in = 12'h101; 
        #20 data_in = 12'h102; 
        #20 data_in = 12'h103; 
        #20 data_in = 12'h104; 
        #20 data_in = 12'h105; 
        #20 data_in = 12'h106; 
        #20 data_in = 12'h107; 
        #20 data_in = 12'h108; 
        #20 data_in = 12'h109; 
        #20 data_in = 12'h10a; 
        #20 data_in = 12'h10b; 
        #20 data_in = 12'h10c; 
        #20 data_in = 12'h10d; 
        #20 data_in = 12'h10e; 
        #20 data_in = 12'h10f; 
        #20 data_in = 12'h110; 
        #20 data_in = 12'h111; 
        #20 data_in = 12'h112; 
        #20 data_in = 12'h113; 
        #20 data_in = 12'h114; 
        #20 data_in = 12'h115; 
        #20 data_in = 12'h116; 
        #20 data_in = 12'h117; 
        #20 data_in = 12'h118; 
        #20 data_in = 12'h119; 
        #20 data_in = 12'h11a; 
        #20 data_in = 12'h11b; 
        #20 data_in = 12'h11c; 
        #20 data_in = 12'h11d; 
        #20 data_in = 12'h11e; 
        #20 data_in = 12'h11f; 
        #20 data_in = 12'h120; 
        #20 data_in = 12'h121; 
        #20 data_in = 12'h122; 
        #20 data_in = 12'h123; 
        #20 data_in = 12'h124; 
        #20 data_in = 12'h125; 
        #20 data_in = 12'h126; 
        #20 data_in = 12'h127; 
        #20 data_in = 12'h128; 
        #20 data_in = 12'h129; 
        #20 data_in = 12'h12a; 
        #20 data_in = 12'h12b; 
        #20 data_in = 12'h12c; 
        #20 data_in = 12'h12d; 
        #20 data_in = 12'h12e; 
        #20 data_in = 12'h12f; 
        #20 data_in = 12'h130; 
        #20 data_in = 12'h131; 
        #20 data_in = 12'h132; 
        #20 data_in = 12'h133; 
        #20 data_in = 12'h134; 
        #20 data_in = 12'h135; 
        #20 data_in = 12'h136; 
        #20 data_in = 12'h137; 
        #20 data_in = 12'h138; 
        #20 data_in = 12'h139; 
        #20 data_in = 12'h13a; 
        #20 data_in = 12'h13b; 
        #20 data_in = 12'h13c; 
        #20 data_in = 12'h13d; 
        #20 data_in = 12'h13e; 
        #20 data_in = 12'h13f; 
        #20 data_in = 12'h140; 
        #20 data_in = 12'h141; 
        #20 data_in = 12'h142; 
        #20 data_in = 12'h143; 
        #20 data_in = 12'h144; 
        #20 data_in = 12'h145; 
        #20 data_in = 12'h146; 
        #20 data_in = 12'h147; 
        #20 data_in = 12'h148; 
        #20 data_in = 12'h149; 
        #20 data_in = 12'h14a; 
        #20 data_in = 12'h14b; 
        #20 data_in = 12'h14c; 
        #20 data_in = 12'h14d; 
        #20 data_in = 12'h14e; 
        #20 data_in = 12'h14f; 
        #20 data_in = 12'h150; 
        #20 data_in = 12'h151; 
        #20 data_in = 12'h152; 
        #20 data_in = 12'h153; 
        #20 data_in = 12'h154; 
        #20 data_in = 12'h155; 
        #20 data_in = 12'h156; 
        #20 data_in = 12'h157; 
        #20 data_in = 12'h158; 
        #20 data_in = 12'h159; 
        #20 data_in = 12'h15a; 
        #20 data_in = 12'h15b; 
        #20 data_in = 12'h15c; 
        #20 data_in = 12'h15d; 
        #20 data_in = 12'h15e; 
        #20 data_in = 12'h15f; 
        #20 data_in = 12'h160; 
        #20 data_in = 12'h161; 
        #20 data_in = 12'h162; 
        #20 data_in = 12'h163; 
        #20 data_in = 12'h164; 
        #20 data_in = 12'h165; 
        #20 data_in = 12'h166; 
        #20 data_in = 12'h167; 
        #20 data_in = 12'h168; 
        #20 data_in = 12'h169; 
        #20 data_in = 12'h16a; 
        #20 data_in = 12'h16b; 
        #20 data_in = 12'h16c; 
        #20 data_in = 12'h16d; 
        #20 data_in = 12'h16e; 
        #20 data_in = 12'h16f; 
        #20 data_in = 12'h170; 
        #20 data_in = 12'h171; 
        #20 data_in = 12'h172; 
        #20 data_in = 12'h173; 
        #20 data_in = 12'h174; 
        #20 data_in = 12'h175; 
        #20 data_in = 12'h176; 
        #20 data_in = 12'h177; 
        #20 data_in = 12'h178; 
        #20 data_in = 12'h179; 
        #20 data_in = 12'h17a; 
        #20 data_in = 12'h17b; 
        #20 data_in = 12'h17c; 
        #20 data_in = 12'h17d; 
        #20 data_in = 12'h17e; 
        #20 data_in = 12'h17f; 
        #20 data_in = 12'h180; 
        #20 data_in = 12'h181; 
        #20 data_in = 12'h182; 
        #20 data_in = 12'h183; 
        #20 data_in = 12'h184; 
        #20 data_in = 12'h185; 
        #20 data_in = 12'h186; 
        #20 data_in = 12'h187; 
        #20 data_in = 12'h188; 
        #20 data_in = 12'h189; 
        #20 data_in = 12'h18a; 
        #20 data_in = 12'h18b; 
        #20 data_in = 12'h18c; 
        #20 data_in = 12'h18d; 
        #20 data_in = 12'h18e; 
        #20 data_in = 12'h18f; 
        #20 data_in = 12'h190; 
        #20 data_in = 12'h191; 
        #20 data_in = 12'h192; 
        #20 data_in = 12'h193; 
        #20 data_in = 12'h194; 
        #20 data_in = 12'h195; 
        #20 data_in = 12'h196; 
        #20 data_in = 12'h197; 
        #20 data_in = 12'h198; 
        #20 data_in = 12'h199; 
        #20 data_in = 12'h19a; 
        #20 data_in = 12'h19b; 
        #20 data_in = 12'h19c; 
        #20 data_in = 12'h19d; 
        #20 data_in = 12'h19e; 
        #20 data_in = 12'h19f; 
        #20 data_in = 12'h1a0; 
        #20 data_in = 12'h1a1; 
        #20 data_in = 12'h1a2; 
        #20 data_in = 12'h1a3; 
        #20 data_in = 12'h1a4; 
        #20 data_in = 12'h1a5; 
        #20 data_in = 12'h1a6; 
        #20 data_in = 12'h1a7; 
        #20 data_in = 12'h1a8; 
        #20 data_in = 12'h1a9; 
        #20 data_in = 12'h1aa; 
        #20 data_in = 12'h1ab; 
        #20 data_in = 12'h1ac; 
        #20 data_in = 12'h1ad; 
        #20 data_in = 12'h1ae; 
        #20 data_in = 12'h1af; 
        #20 data_in = 12'h1b0; 
        #20 data_in = 12'h1b1; 
        #20 data_in = 12'h1b2; 
        #20 data_in = 12'h1b3; 
        #20 data_in = 12'h1b4; 
        #20 data_in = 12'h1b5; 
        #20 data_in = 12'h1b6; 
        #20 data_in = 12'h1b7; 
        #20 data_in = 12'h1b8; 
        #20 data_in = 12'h1b9; 
        #20 data_in = 12'h1ba; 
        #20 data_in = 12'h1bb; 
        #20 data_in = 12'h1bc; 
        #20 data_in = 12'h1bd; 
        #20 data_in = 12'h1be; 
        #20 data_in = 12'h1bf; 
        #20 data_in = 12'h1c0; 
        #20 data_in = 12'h1c1; 
        #20 data_in = 12'h1c2; 
        #20 data_in = 12'h1c3; 
        #20 data_in = 12'h1c4; 
        #20 data_in = 12'h1c5; 
        #20 data_in = 12'h1c6; 
        #20 data_in = 12'h1c7; 
        #20 data_in = 12'h1c8; 
        #20 data_in = 12'h1c9; 
        #20 data_in = 12'h1ca; 
        #20 data_in = 12'h1cb; 
        #20 data_in = 12'h1cc; 
        #20 data_in = 12'h1cd; 
        #20 data_in = 12'h1ce; 
        #20 data_in = 12'h1cf; 
        #20 data_in = 12'h1d0; 
        #20 data_in = 12'h1d1; 
        #20 data_in = 12'h1d2; 
        #20 data_in = 12'h1d3; 
        #20 data_in = 12'h1d4; 
        #20 data_in = 12'h1d5; 
        #20 data_in = 12'h1d6; 
        #20 data_in = 12'h1d7; 
        #20 data_in = 12'h1d8; 
        #20 data_in = 12'h1d9; 
        #20 data_in = 12'h1da; 
        #20 data_in = 12'h1db; 
        #20 data_in = 12'h1dc; 
        #20 data_in = 12'h1dd; 
        #20 data_in = 12'h1de; 
        #20 data_in = 12'h1df; 
        #20 data_in = 12'h1e0; 
        #20 data_in = 12'h1e1; 
        #20 data_in = 12'h1e2; 
        #20 data_in = 12'h1e3; 
        #20 data_in = 12'h1e4; 
        #20 data_in = 12'h1e5; 
        #20 data_in = 12'h1e6; 
        #20 data_in = 12'h1e7; 
        #20 data_in = 12'h1e8; 
        #20 data_in = 12'h1e9; 
        #20 data_in = 12'h1ea; 
        #20 data_in = 12'h1eb; 
        #20 data_in = 12'h1ec; 
        #20 data_in = 12'h1ed; 
        #20 data_in = 12'h1ee; 
        #20 data_in = 12'h1ef; 
        #20 data_in = 12'h1f0; 
        #20 data_in = 12'h1f1; 
        #20 data_in = 12'h1f2; 
        #20 data_in = 12'h1f3; 
        #20 data_in = 12'h1f4; 
        #20 data_in = 12'h1f5; 
        #20 data_in = 12'h1f6; 
        #20 data_in = 12'h1f7; 
        #20 data_in = 12'h1f8; 
        #20 data_in = 12'h1f9; 
        #20 data_in = 12'h1fa; 
        #20 data_in = 12'h1fb; 
        #20 data_in = 12'h1fc; 
        #20 data_in = 12'h1fd; 
        #20 data_in = 12'h1fe; 
        #20 data_in = 12'h1ff; 
        #20 data_in = 12'h200; 
        #20 data_in = 12'h201; 
        #20 data_in = 12'h202; 
        #20 data_in = 12'h203; 
        #20 data_in = 12'h204; 
        #20 data_in = 12'h205; 
        #20 data_in = 12'h206; 
        #20 data_in = 12'h207; 
        #20 data_in = 12'h208; 
        #20 data_in = 12'h209; 
        #20 data_in = 12'h20a; 
        #20 data_in = 12'h20b; 
        #20 data_in = 12'h20c; 
        #20 data_in = 12'h20d; 
        #20 data_in = 12'h20e; 
        #20 data_in = 12'h20f; 
        #20 data_in = 12'h210; 
        #20 data_in = 12'h211; 
        #20 data_in = 12'h212; 
        #20 data_in = 12'h213; 
        #20 data_in = 12'h214; 
        #20 data_in = 12'h215; 
        #20 data_in = 12'h216; 
        #20 data_in = 12'h217; 
        #20 data_in = 12'h218; 
        #20 data_in = 12'h219; 
        #20 data_in = 12'h21a; 
        #20 data_in = 12'h21b; 
        #20 data_in = 12'h21c; 
        #20 data_in = 12'h21d; 
        #20 data_in = 12'h21e; 
        #20 data_in = 12'h21f; 
        #20 data_in = 12'h220; 
        #20 data_in = 12'h221; 
        #20 data_in = 12'h222; 
        #20 data_in = 12'h223; 
        #20 data_in = 12'h224; 
        #20 data_in = 12'h225; 
        #20 data_in = 12'h226; 
        #20 data_in = 12'h227; 
        #20 data_in = 12'h228; 
        #20 data_in = 12'h229; 
        #20 data_in = 12'h22a; 
        #20 data_in = 12'h22b; 
        #20 data_in = 12'h22c; 
        #20 data_in = 12'h22d; 
        #20 data_in = 12'h22e; 
        #20 data_in = 12'h22f; 
        #20 data_in = 12'h230; 
        #20 data_in = 12'h231; 
        #20 data_in = 12'h232; 
        #20 data_in = 12'h233; 
        #20 data_in = 12'h234; 
        #20 data_in = 12'h235; 
        #20 data_in = 12'h236; 
        #20 data_in = 12'h237; 
        #20 data_in = 12'h238; 
        #20 data_in = 12'h239; 
        #20 data_in = 12'h23a; 
        #20 data_in = 12'h23b; 
        #20 data_in = 12'h23c; 
        #20 data_in = 12'h23d; 
        #20 data_in = 12'h23e; 
        #20 data_in = 12'h23f; 
        #20 data_in = 12'h240; 
        #20 data_in = 12'h241; 
        #20 data_in = 12'h242; 
        #20 data_in = 12'h243; 
        #20 data_in = 12'h244; 
        #20 data_in = 12'h245; 
        #20 data_in = 12'h246; 
        #20 data_in = 12'h247; 
        #20 data_in = 12'h248; 
        #20 data_in = 12'h249; 
        #20 data_in = 12'h24a; 
        #20 data_in = 12'h24b; 
        #20 data_in = 12'h24c; 
        #20 data_in = 12'h24d; 
        #20 data_in = 12'h24e; 
        #20 data_in = 12'h24f; 
        #20 data_in = 12'h250; 
        #20 data_in = 12'h251; 
        #20 data_in = 12'h252; 
        #20 data_in = 12'h253; 
        #20 data_in = 12'h254; 
        #20 data_in = 12'h255; 
        #20 data_in = 12'h256; 
        #20 data_in = 12'h257; 
        #20 data_in = 12'h258; 
        #20 data_in = 12'h259; 
        #20 data_in = 12'h25a; 
        #20 data_in = 12'h25b; 
        #20 data_in = 12'h25c; 
        #20 data_in = 12'h25d; 
        #20 data_in = 12'h25e; 
        #20 data_in = 12'h25f; 
        #20 data_in = 12'h260; 
        #20 data_in = 12'h261; 
        #20 data_in = 12'h262; 
        #20 data_in = 12'h263; 
        #20 data_in = 12'h264; 
        #20 data_in = 12'h265; 
        #20 data_in = 12'h266; 
        #20 data_in = 12'h267; 
        #20 data_in = 12'h268; 
        #20 data_in = 12'h269; 
        #20 data_in = 12'h26a; 
        #20 data_in = 12'h26b; 
        #20 data_in = 12'h26c; 
        #20 data_in = 12'h26d; 
        #20 data_in = 12'h26e; 
        #20 data_in = 12'h26f; 
        #20 data_in = 12'h270; 
        #20 data_in = 12'h271; 
        #20 data_in = 12'h272; 
        #20 data_in = 12'h273; 
        #20 data_in = 12'h274; 
        #20 data_in = 12'h275; 
        #20 data_in = 12'h276; 
        #20 data_in = 12'h277; 
        #20 data_in = 12'h278; 
        #20 data_in = 12'h279; 
        #20 data_in = 12'h27a; 
        #20 data_in = 12'h27b; 
        #20 data_in = 12'h27c; 
        #20 data_in = 12'h27d; 
        #20 data_in = 12'h27e; 
        #20 data_in = 12'h27f; 
        #20 data_in = 12'h280; 
        #20 data_in = 12'h281; 
        #20 data_in = 12'h282; 
        #20 data_in = 12'h283; 
        #20 data_in = 12'h284; 
        #20 data_in = 12'h285; 
        #20 data_in = 12'h286; 
        #20 data_in = 12'h287; 
        #20 data_in = 12'h288; 
        #20 data_in = 12'h289; 
        #20 data_in = 12'h28a; 
        #20 data_in = 12'h28b; 
        #20 data_in = 12'h28c; 
        #20 data_in = 12'h28d; 
        #20 data_in = 12'h28e; 
        #20 data_in = 12'h28f; 
        #20 data_in = 12'h290; 
        #20 data_in = 12'h291; 
        #20 data_in = 12'h292; 
        #20 data_in = 12'h293; 
        #20 data_in = 12'h294; 
        #20 data_in = 12'h295; 
        #20 data_in = 12'h296; 
        #20 data_in = 12'h297; 
        #20 data_in = 12'h298; 
        #20 data_in = 12'h299; 
        #20 data_in = 12'h29a; 
        #20 data_in = 12'h29b; 
        #20 data_in = 12'h29c; 
        #20 data_in = 12'h29d; 
        #20 data_in = 12'h29e; 
        #20 data_in = 12'h29f; 
        #20 data_in = 12'h2a0; 
        #20 data_in = 12'h2a1; 
        #20 data_in = 12'h2a2; 
        #20 data_in = 12'h2a3; 
        #20 data_in = 12'h2a4; 
        #20 data_in = 12'h2a5; 
        #20 data_in = 12'h2a6; 
        #20 data_in = 12'h2a7; 
        #20 data_in = 12'h2a8; 
        #20 data_in = 12'h2a9; 
        #20 data_in = 12'h2aa; 
        #20 data_in = 12'h2ab; 
        #20 data_in = 12'h2ac; 
        #20 data_in = 12'h2ad; 
        #20 data_in = 12'h2ae; 
        #20 data_in = 12'h2af; 
        #20 data_in = 12'h2b0; 
        #20 data_in = 12'h2b1; 
        #20 data_in = 12'h2b2; 
        #20 data_in = 12'h2b3; 
        #20 data_in = 12'h2b4; 
        #20 data_in = 12'h2b5; 
        #20 data_in = 12'h2b6; 
        #20 data_in = 12'h2b7; 
        #20 data_in = 12'h2b8; 
        #20 data_in = 12'h2b9; 
        #20 data_in = 12'h2ba; 
        #20 data_in = 12'h2bb; 
        #20 data_in = 12'h2bc; 
        #20 data_in = 12'h2bd; 
        #20 data_in = 12'h2be; 
        #20 data_in = 12'h2bf; 
        #20 data_in = 12'h2c0; 
        #20 data_in = 12'h2c1; 
        #20 data_in = 12'h2c2; 
        #20 data_in = 12'h2c3; 
        #20 data_in = 12'h2c4; 
        #20 data_in = 12'h2c5; 
        #20 data_in = 12'h2c6; 
        #20 data_in = 12'h2c7; 
        #20 data_in = 12'h2c8; 
        #20 data_in = 12'h2c9; 
        #20 data_in = 12'h2ca; 
        #20 data_in = 12'h2cb; 
        #20 data_in = 12'h2cc; 
        #20 data_in = 12'h2cd; 
        #20 data_in = 12'h2ce; 
        #20 data_in = 12'h2cf; 
        #20 data_in = 12'h2d0; 
        #20 data_in = 12'h2d1; 
        #20 data_in = 12'h2d2; 
        #20 data_in = 12'h2d3; 
        #20 data_in = 12'h2d4; 
        #20 data_in = 12'h2d5; 
        #20 data_in = 12'h2d6; 
        #20 data_in = 12'h2d7; 
        #20 data_in = 12'h2d8; 
        #20 data_in = 12'h2d9; 
        #20 data_in = 12'h2da; 
        #20 data_in = 12'h2db; 
        #20 data_in = 12'h2dc; 
        #20 data_in = 12'h2dd; 
        #20 data_in = 12'h2de; 
        #20 data_in = 12'h2df; 
        #20 data_in = 12'h2e0; 
        #20 data_in = 12'h2e1; 
        #20 data_in = 12'h2e2; 
        #20 data_in = 12'h2e3; 
        #20 data_in = 12'h2e4; 
        #20 data_in = 12'h2e5; 
        #20 data_in = 12'h2e6; 
        #20 data_in = 12'h2e7; 
        #20 data_in = 12'h2e8; 
        #20 data_in = 12'h2e9; 
        #20 data_in = 12'h2ea; 
        #20 data_in = 12'h2eb; 
        #20 data_in = 12'h2ec; 
        #20 data_in = 12'h2ed; 
        #20 data_in = 12'h2ee; 
        #20 data_in = 12'h2ef; 
        #20 data_in = 12'h2f0; 
        #20 data_in = 12'h2f1; 
        #20 data_in = 12'h2f2; 
        #20 data_in = 12'h2f3; 
        #20 data_in = 12'h2f4; 
        #20 data_in = 12'h2f5; 
        #20 data_in = 12'h2f6; 
        #20 data_in = 12'h2f7; 
        #20 data_in = 12'h2f8; 
        #20 data_in = 12'h2f9; 
        #20 data_in = 12'h2fa; 
        #20 data_in = 12'h2fb; 
        #20 data_in = 12'h2fc; 
        #20 data_in = 12'h2fd; 
        #20 data_in = 12'h2fe; 
        #20 data_in = 12'h2ff; 
        #20 data_in = 12'h300; 
        #20 data_in = 12'h301; 
        #20 data_in = 12'h302; 
        #20 data_in = 12'h303; 
        #20 data_in = 12'h304; 
        #20 data_in = 12'h305; 
        #20 data_in = 12'h306; 
        #20 data_in = 12'h307; 
        #20 data_in = 12'h308; 
        #20 data_in = 12'h309; 
        #20 data_in = 12'h30a; 
        #20 data_in = 12'h30b; 
        #20 data_in = 12'h30c; 
        #20 data_in = 12'h30d; 
        #20 data_in = 12'h30e; 
        #20 data_in = 12'h30f; 
        #20 data_in = 12'h310; 
        #20 data_in = 12'h311; 
        #20 data_in = 12'h312; 
        #20 data_in = 12'h313; 
        #20 data_in = 12'h314; 
        #20 data_in = 12'h315; 
        #20 data_in = 12'h316; 
        #20 data_in = 12'h317; 
        #20 data_in = 12'h318; 
        #20 data_in = 12'h319; 
        #20 data_in = 12'h31a; 
        #20 data_in = 12'h31b; 
        #20 data_in = 12'h31c; 
        #20 data_in = 12'h31d; 
        #20 data_in = 12'h31e; 
        #20 data_in = 12'h31f; 
        #20 data_in = 12'h320; 
        #20 data_in = 12'h321; 
        #20 data_in = 12'h322; 
        #20 data_in = 12'h323; 
        #20 data_in = 12'h324; 
        #20 data_in = 12'h325; 
        #20 data_in = 12'h326; 
        #20 data_in = 12'h327; 
        #20 data_in = 12'h328; 
        #20 data_in = 12'h329; 
        #20 data_in = 12'h32a; 
        #20 data_in = 12'h32b; 
        #20 data_in = 12'h32c; 
        #20 data_in = 12'h32d; 
        #20 data_in = 12'h32e; 
        #20 data_in = 12'h32f; 
        #20 data_in = 12'h330; 
        #20 data_in = 12'h331; 
        #20 data_in = 12'h332; 
        #20 data_in = 12'h333; 
        #20 data_in = 12'h334; 
        #20 data_in = 12'h335; 
        #20 data_in = 12'h336; 
        #20 data_in = 12'h337; 
        #20 data_in = 12'h338; 
        #20 data_in = 12'h339; 
        #20 data_in = 12'h33a; 
        #20 data_in = 12'h33b; 
        #20 data_in = 12'h33c; 
        #20 data_in = 12'h33d; 
        #20 data_in = 12'h33e; 
        #20 data_in = 12'h33f; 
        #20 data_in = 12'h340; 
        #20 data_in = 12'h341; 
        #20 data_in = 12'h342; 
        #20 data_in = 12'h343; 
        #20 data_in = 12'h344; 
        #20 data_in = 12'h345; 
        #20 data_in = 12'h346; 
        #20 data_in = 12'h347; 
        #20 data_in = 12'h348; 
        #20 data_in = 12'h349; 
        #20 data_in = 12'h34a; 
        #20 data_in = 12'h34b; 
        #20 data_in = 12'h34c; 
        #20 data_in = 12'h34d; 
        #20 data_in = 12'h34e; 
        #20 data_in = 12'h34f; 
        #20 data_in = 12'h350; 
        #20 data_in = 12'h351; 
        #20 data_in = 12'h352; 
        #20 data_in = 12'h353; 
        #20 data_in = 12'h354; 
        #20 data_in = 12'h355; 
        #20 data_in = 12'h356; 
        #20 data_in = 12'h357; 
        #20 data_in = 12'h358; 
        #20 data_in = 12'h359; 
        #20 data_in = 12'h35a; 
        #20 data_in = 12'h35b; 
        #20 data_in = 12'h35c; 
        #20 data_in = 12'h35d; 
        #20 data_in = 12'h35e; 
        #20 data_in = 12'h35f; 
        #20 data_in = 12'h360; 
        #20 data_in = 12'h361; 
        #20 data_in = 12'h362; 
        #20 data_in = 12'h363; 
        #20 data_in = 12'h364; 
        #20 data_in = 12'h365; 
        #20 data_in = 12'h366; 
        #20 data_in = 12'h367; 
        #20 data_in = 12'h368; 
        #20 data_in = 12'h369; 
        #20 data_in = 12'h36a; 
        #20 data_in = 12'h36b; 
        #20 data_in = 12'h36c; 
        #20 data_in = 12'h36d; 
        #20 data_in = 12'h36e; 
        #20 data_in = 12'h36f; 
        #20 data_in = 12'h370; 
        #20 data_in = 12'h371; 
        #20 data_in = 12'h372; 
        #20 data_in = 12'h373; 
        #20 data_in = 12'h374; 
        #20 data_in = 12'h375; 
        #20 data_in = 12'h376; 
        #20 data_in = 12'h377; 
        #20 data_in = 12'h378; 
        #20 data_in = 12'h379; 
        #20 data_in = 12'h37a; 
        #20 data_in = 12'h37b; 
        #20 data_in = 12'h37c; 
        #20 data_in = 12'h37d; 
        #20 data_in = 12'h37e; 
        #20 data_in = 12'h37f; 
        #20 data_in = 12'h380; 
        #20 data_in = 12'h381; 
        #20 data_in = 12'h382; 
        #20 data_in = 12'h383; 
        #20 data_in = 12'h384; 
        #20 data_in = 12'h385; 
        #20 data_in = 12'h386; 
        #20 data_in = 12'h387; 
        #20 data_in = 12'h388; 
        #20 data_in = 12'h389; 
        #20 data_in = 12'h38a; 
        #20 data_in = 12'h38b; 
        #20 data_in = 12'h38c; 
        #20 data_in = 12'h38d; 
        #20 data_in = 12'h38e; 
        #20 data_in = 12'h38f; 
        #20 data_in = 12'h390; 
        #20 data_in = 12'h391; 
        #20 data_in = 12'h392; 
        #20 data_in = 12'h393; 
        #20 data_in = 12'h394; 
        #20 data_in = 12'h395; 
        #20 data_in = 12'h396; 
        #20 data_in = 12'h397; 
        #20 data_in = 12'h398; 
        #20 data_in = 12'h399; 
        #20 data_in = 12'h39a; 
        #20 data_in = 12'h39b; 
        #20 data_in = 12'h39c; 
        #20 data_in = 12'h39d; 
        #20 data_in = 12'h39e; 
        #20 data_in = 12'h39f; 
        #20 data_in = 12'h3a0; 
        #20 data_in = 12'h3a1; 
        #20 data_in = 12'h3a2; 
        #20 data_in = 12'h3a3; 
        #20 data_in = 12'h3a4; 
        #20 data_in = 12'h3a5; 
        #20 data_in = 12'h3a6; 
        #20 data_in = 12'h3a7; 
        #20 data_in = 12'h3a8; 
        #20 data_in = 12'h3a9; 
        #20 data_in = 12'h3aa; 
        #20 data_in = 12'h3ab; 
        #20 data_in = 12'h3ac; 
        #20 data_in = 12'h3ad; 
        #20 data_in = 12'h3ae; 
        #20 data_in = 12'h3af; 
        #20 data_in = 12'h3b0; 
        #20 data_in = 12'h3b1; 
        #20 data_in = 12'h3b2; 
        #20 data_in = 12'h3b3; 
        #20 data_in = 12'h3b4; 
        #20 data_in = 12'h3b5; 
        #20 data_in = 12'h3b6; 
        #20 data_in = 12'h3b7; 
        #20 data_in = 12'h3b8; 
        #20 data_in = 12'h3b9; 
        #20 data_in = 12'h3ba; 
        #20 data_in = 12'h3bb; 
        #20 data_in = 12'h3bc; 
        #20 data_in = 12'h3bd; 
        #20 data_in = 12'h3be; 
        #20 data_in = 12'h3bf; 
        #20 data_in = 12'h3c0; 
        #20 data_in = 12'h3c1; 
        #20 data_in = 12'h3c2; 
        #20 data_in = 12'h3c3; 
        #20 data_in = 12'h3c4; 
        #20 data_in = 12'h3c5; 
        #20 data_in = 12'h3c6; 
        #20 data_in = 12'h3c7; 
        #20 data_in = 12'h3c8; 
        #20 data_in = 12'h3c9; 
        #20 data_in = 12'h3ca; 
        #20 data_in = 12'h3cb; 
        #20 data_in = 12'h3cc; 
        #20 data_in = 12'h3cd; 
        #20 data_in = 12'h3ce; 
        #20 data_in = 12'h3cf; 
        #20 data_in = 12'h3d0; 
        #20 data_in = 12'h3d1; 
        #20 data_in = 12'h3d2; 
        #20 data_in = 12'h3d3; 
        #20 data_in = 12'h3d4; 
        #20 data_in = 12'h3d5; 
        #20 data_in = 12'h3d6; 
        #20 data_in = 12'h3d7; 
        #20 data_in = 12'h3d8; 
        #20 data_in = 12'h3d9; 
        #20 data_in = 12'h3da; 
        #20 data_in = 12'h3db; 
        #20 data_in = 12'h3dc; 
        #20 data_in = 12'h3dd; 
        #20 data_in = 12'h3de; 
        #20 data_in = 12'h3df; 
        #20 data_in = 12'h3e0; 
        #20 data_in = 12'h3e1; 
        #20 data_in = 12'h3e2; 
        #20 data_in = 12'h3e3; 
        #20 data_in = 12'h3e4; 
        #20 data_in = 12'h3e5; 
        #20 data_in = 12'h3e6; 
        #20 data_in = 12'h3e7; 
        #20 data_in = 12'h3e8; 
        #20 data_in = 12'h3e9; 
        #20 data_in = 12'h3ea; 
        #20 data_in = 12'h3eb; 
        #20 data_in = 12'h3ec; 
        #20 data_in = 12'h3ed; 
        #20 data_in = 12'h3ee; 
        #20 data_in = 12'h3ef; 
        #20 data_in = 12'h3f0; 
        #20 data_in = 12'h3f1; 
        #20 data_in = 12'h3f2; 
        #20 data_in = 12'h3f3; 
        #20 data_in = 12'h3f4; 
        #20 data_in = 12'h3f5; 
        #20 data_in = 12'h3f6; 
        #20 data_in = 12'h3f7; 
        #20 data_in = 12'h3f8; 
        #20 data_in = 12'h3f9; 
        #20 data_in = 12'h3fa; 
        #20 data_in = 12'h3fb; 
        #20 data_in = 12'h3fc; 
        #20 data_in = 12'h3fd; 
        #20 data_in = 12'h3fe; 
        #20 data_in = 12'h3ff;		
        #20 data_in = 12'h400; 
        #20 data_in = 12'h401;
        #20 data_in = 12'h402; 
        #20 data_in = 12'h403; 
        #20 data_in = 12'h404;
        #20 data_in = 12'h405; 
        #20 data_in = 12'h406;
        #20 data_in = 12'h407; 
        #20 data_in = 12'h408; 
        #20 data_in = 12'h409; 
        #20 data_in = 12'h40a; 
        #20 data_in = 12'h40b; 
        #20 data_in = 12'h40c; 
        #20 data_in = 12'h40d; 
        #20 data_in = 12'h40e; 
        #20 data_in = 12'h40f; 
        #20 data_in = 12'h410; 
        #20 data_in = 12'h411; 
        #20 data_in = 12'h412; 
        #20 data_in = 12'h413; 
        #20 data_in = 12'h414; 
        #20 data_in = 12'h415; 
        #20 data_in = 12'h416; 
        #20 data_in = 12'h417; 
        #20 data_in = 12'h418; 
        #20 data_in = 12'h419; 
        #20 data_in = 12'h41a; 
        #20 data_in = 12'h41b; 
        #20 data_in = 12'h41c; 
        #20 data_in = 12'h41d; 
        #20 data_in = 12'h41e; 
        #20 data_in = 12'h41f; 
        #20 data_in = 12'h420; 
        #20 data_in = 12'h421; 
        #20 data_in = 12'h422; 
        #20 data_in = 12'h423; 
        #20 data_in = 12'h424; 
        #20 data_in = 12'h425; 
        #20 data_in = 12'h426; 
        #20 data_in = 12'h427; 
        #20 data_in = 12'h428; 
        #20 data_in = 12'h429; 
        #20 data_in = 12'h42a; 
        #20 data_in = 12'h42b; 
        #20 data_in = 12'h42c; 
        #20 data_in = 12'h42d; 
        #20 data_in = 12'h42e; 
        #20 data_in = 12'h42f; 
        #20 data_in = 12'h430; 
        #20 data_in = 12'h431; 
        #20 data_in = 12'h432; 
        #20 data_in = 12'h433; 
        #20 data_in = 12'h434; 
        #20 data_in = 12'h435; 
        #20 data_in = 12'h436; 
        #20 data_in = 12'h437; 
        #20 data_in = 12'h438; 
        #20 data_in = 12'h439; 
        #20 data_in = 12'h43a; 
        #20 data_in = 12'h43b; 
        #20 data_in = 12'h43c; 
        #20 data_in = 12'h43d; 
        #20 data_in = 12'h43e; 
        #20 data_in = 12'h43f; 
        #20 data_in = 12'h440; 
        #20 data_in = 12'h441; 
        #20 data_in = 12'h442; 
        #20 data_in = 12'h443; 
        #20 data_in = 12'h444; 
        #20 data_in = 12'h445; 
        #20 data_in = 12'h446; 
        #20 data_in = 12'h447; 
        #20 data_in = 12'h448; 
        #20 data_in = 12'h449; 
        #20 data_in = 12'h44a; 
        #20 data_in = 12'h44b; 
        #20 data_in = 12'h44c; 
        #20 data_in = 12'h44d; 
        #20 data_in = 12'h44e; 
        #20 data_in = 12'h44f; 
        #20 data_in = 12'h450; 
        #20 data_in = 12'h451; 
        #20 data_in = 12'h452; 
        #20 data_in = 12'h453; 
        #20 data_in = 12'h454; 
        #20 data_in = 12'h455; 
        #20 data_in = 12'h456; 
        #20 data_in = 12'h457; 
        #20 data_in = 12'h458; 
        #20 data_in = 12'h459; 
        #20 data_in = 12'h45a; 
        #20 data_in = 12'h45b; 
        #20 data_in = 12'h45c; 
        #20 data_in = 12'h45d; 
        #20 data_in = 12'h45e; 
        #20 data_in = 12'h45f; 
        #20 data_in = 12'h460; 
        #20 data_in = 12'h461; 
        #20 data_in = 12'h462; 
        #20 data_in = 12'h463; 
        #20 data_in = 12'h464; 
        #20 data_in = 12'h465; 
        #20 data_in = 12'h466; 
        #20 data_in = 12'h467; 
        #20 data_in = 12'h468; 
        #20 data_in = 12'h469; 
        #20 data_in = 12'h46a; 
        #20 data_in = 12'h46b; 
        #20 data_in = 12'h46c; 
        #20 data_in = 12'h46d; 
        #20 data_in = 12'h46e; 
        #20 data_in = 12'h46f; 
        #20 data_in = 12'h470; 
        #20 data_in = 12'h471; 
        #20 data_in = 12'h472; 
        #20 data_in = 12'h473; 
        #20 data_in = 12'h474; 
        #20 data_in = 12'h475; 
        #20 data_in = 12'h476; 
        #20 data_in = 12'h477; 
        #20 data_in = 12'h478; 
        #20 data_in = 12'h479; 
        #20 data_in = 12'h47a; 
        #20 data_in = 12'h47b; 
        #20 data_in = 12'h47c; 
        #20 data_in = 12'h47d; 
        #20 data_in = 12'h47e; 
        #20 data_in = 12'h47f; 
        #20 data_in = 12'h480; 
        #20 data_in = 12'h481; 
        #20 data_in = 12'h482; 
        #20 data_in = 12'h483; 
        #20 data_in = 12'h484; 
        #20 data_in = 12'h485; 
        #20 data_in = 12'h486; 
        #20 data_in = 12'h487; 
        #20 data_in = 12'h488; 
        #20 data_in = 12'h489; 
        #20 data_in = 12'h48a; 
        #20 data_in = 12'h48b; 
        #20 data_in = 12'h48c; 
        #20 data_in = 12'h48d; 
        #20 data_in = 12'h48e; 
        #20 data_in = 12'h48f; 
        #20 data_in = 12'h490; 
        #20 data_in = 12'h491; 
        #20 data_in = 12'h492; 
        #20 data_in = 12'h493; 
        #20 data_in = 12'h494; 
        #20 data_in = 12'h495; 
        #20 data_in = 12'h496; 
        #20 data_in = 12'h497; 
        #20 data_in = 12'h498; 
        #20 data_in = 12'h499; 
        #20 data_in = 12'h49a; 
        #20 data_in = 12'h49b; 
        #20 data_in = 12'h49c; 
        #20 data_in = 12'h49d; 
        #20 data_in = 12'h49e; 
        #20 data_in = 12'h49f; 
        #20 data_in = 12'h4a0; 
        #20 data_in = 12'h4a1; 
        #20 data_in = 12'h4a2; 
        #20 data_in = 12'h4a3; 
        #20 data_in = 12'h4a4; 
        #20 data_in = 12'h4a5; 
        #20 data_in = 12'h4a6; 
        #20 data_in = 12'h4a7; 
        #20 data_in = 12'h4a8; 
        #20 data_in = 12'h4a9; 
        #20 data_in = 12'h4aa; 
        #20 data_in = 12'h4ab; 
        #20 data_in = 12'h4ac; 
        #20 data_in = 12'h4ad; 
        #20 data_in = 12'h4ae; 
        #20 data_in = 12'h4af; 
        #20 data_in = 12'h4b0; 
        #20 data_in = 12'h4b1; 
        #20 data_in = 12'h4b2; 
        #20 data_in = 12'h4b3; 
        #20 data_in = 12'h4b4; 
        #20 data_in = 12'h4b5; 
        #20 data_in = 12'h4b6; 
        #20 data_in = 12'h4b7; 
        #20 data_in = 12'h4b8; 
        #20 data_in = 12'h4b9; 
        #20 data_in = 12'h4ba; 
        #20 data_in = 12'h4bb; 
        #20 data_in = 12'h4bc; 
        #20 data_in = 12'h4bd; 
        #20 data_in = 12'h4be; 
        #20 data_in = 12'h4bf; 
        #20 data_in = 12'h4c0; 
        #20 data_in = 12'h4c1; 
        #20 data_in = 12'h4c2; 
        #20 data_in = 12'h4c3; 
        #20 data_in = 12'h4c4; 
        #20 data_in = 12'h4c5; 
        #20 data_in = 12'h4c6; 
        #20 data_in = 12'h4c7; 
        #20 data_in = 12'h4c8; 
        #20 data_in = 12'h4c9; 
        #20 data_in = 12'h4ca; 
        #20 data_in = 12'h4cb; 
        #20 data_in = 12'h4cc; 
        #20 data_in = 12'h4cd; 
        #20 data_in = 12'h4ce; 
        #20 data_in = 12'h4cf; 
        #20 data_in = 12'h4d0; 
        #20 data_in = 12'h4d1; 
        #20 data_in = 12'h4d2; 
        #20 data_in = 12'h4d3; 
        #20 data_in = 12'h4d4; 
        #20 data_in = 12'h4d5; 
        #20 data_in = 12'h4d6; 
        #20 data_in = 12'h4d7; 
        #20 data_in = 12'h4d8; 
        #20 data_in = 12'h4d9; 
        #20 data_in = 12'h4da; 
        #20 data_in = 12'h4db; 
        #20 data_in = 12'h4dc; 
        #20 data_in = 12'h4dd; 
        #20 data_in = 12'h4de; 
        #20 data_in = 12'h4df; 
        #20 data_in = 12'h4e0; 
        #20 data_in = 12'h4e1; 
        #20 data_in = 12'h4e2; 
        #20 data_in = 12'h4e3; 
        #20 data_in = 12'h4e4; 
        #20 data_in = 12'h4e5; 
        #20 data_in = 12'h4e6; 
        #20 data_in = 12'h4e7; 
        #20 data_in = 12'h4e8; 
        #20 data_in = 12'h4e9; 
        #20 data_in = 12'h4ea; 
        #20 data_in = 12'h4eb; 
        #20 data_in = 12'h4ec; 
        #20 data_in = 12'h4ed; 
        #20 data_in = 12'h4ee; 
        #20 data_in = 12'h4ef; 
        #20 data_in = 12'h4f0; 
        #20 data_in = 12'h4f1; 
        #20 data_in = 12'h4f2; 
        #20 data_in = 12'h4f3; 
        #20 data_in = 12'h4f4; 
        #20 data_in = 12'h4f5; 
        #20 data_in = 12'h4f6; 
        #20 data_in = 12'h4f7; 
        #20 data_in = 12'h4f8; 
        #20 data_in = 12'h4f9; 
        #20 data_in = 12'h4fa; 
        #20 data_in = 12'h4fb; 
        #20 data_in = 12'h4fc; 
        #20 data_in = 12'h4fd; 
        #20 data_in = 12'h4fe; 
        #20 data_in = 12'h4ff; 
        #20 data_in = 12'h500; 
        #20 data_in = 12'h501; 
        #20 data_in = 12'h502; 
        #20 data_in = 12'h503; 
        #20 data_in = 12'h504; 
        #20 data_in = 12'h505; 
        #20 data_in = 12'h506; 
        #20 data_in = 12'h507; 
        #20 data_in = 12'h508; 
        #20 data_in = 12'h509; 
        #20 data_in = 12'h50a; 
        #20 data_in = 12'h50b; 
        #20 data_in = 12'h50c; 
        #20 data_in = 12'h50d; 
        #20 data_in = 12'h50e; 
        #20 data_in = 12'h50f; 
        #20 data_in = 12'h510; 
        #20 data_in = 12'h511; 
        #20 data_in = 12'h512; 
        #20 data_in = 12'h513; 
        #20 data_in = 12'h514; 
        #20 data_in = 12'h515; 
        #20 data_in = 12'h516; 
        #20 data_in = 12'h517; 
        #20 data_in = 12'h518; 
        #20 data_in = 12'h519; 
        #20 data_in = 12'h51a; 
        #20 data_in = 12'h51b; 
        #20 data_in = 12'h51c; 
        #20 data_in = 12'h51d; 
        #20 data_in = 12'h51e; 
        #20 data_in = 12'h51f; 
        #20 data_in = 12'h520; 
        #20 data_in = 12'h521; 
        #20 data_in = 12'h522; 
        #20 data_in = 12'h523; 
        #20 data_in = 12'h524; 
        #20 data_in = 12'h525; 
        #20 data_in = 12'h526; 
        #20 data_in = 12'h527; 
        #20 data_in = 12'h528; 
        #20 data_in = 12'h529; 
        #20 data_in = 12'h52a; 
        #20 data_in = 12'h52b; 
        #20 data_in = 12'h52c; 
        #20 data_in = 12'h52d; 
        #20 data_in = 12'h52e; 
        #20 data_in = 12'h52f; 
        #20 data_in = 12'h530; 
        #20 data_in = 12'h531; 
        #20 data_in = 12'h532; 
        #20 data_in = 12'h533; 
        #20 data_in = 12'h534; 
        #20 data_in = 12'h535; 
        #20 data_in = 12'h536; 
        #20 data_in = 12'h537; 
        #20 data_in = 12'h538; 
        #20 data_in = 12'h539; 
        #20 data_in = 12'h53a; 
        #20 data_in = 12'h53b; 
        #20 data_in = 12'h53c; 
        #20 data_in = 12'h53d; 
        #20 data_in = 12'h53e; 
        #20 data_in = 12'h53f; 
        #20 data_in = 12'h540; 
        #20 data_in = 12'h541; 
        #20 data_in = 12'h542; 
        #20 data_in = 12'h543; 
        #20 data_in = 12'h544; 
        #20 data_in = 12'h545; 
        #20 data_in = 12'h546; 
        #20 data_in = 12'h547; 
        #20 data_in = 12'h548; 
        #20 data_in = 12'h549; 
        #20 data_in = 12'h54a; 
        #20 data_in = 12'h54b; 
        #20 data_in = 12'h54c; 
        #20 data_in = 12'h54d; 
        #20 data_in = 12'h54e; 
        #20 data_in = 12'h54f; 
        #20 data_in = 12'h550; 
        #20 data_in = 12'h551; 
        #20 data_in = 12'h552; 
        #20 data_in = 12'h553; 
        #20 data_in = 12'h554; 
        #20 data_in = 12'h555; 
        #20 data_in = 12'h556; 
        #20 data_in = 12'h557; 
        #20 data_in = 12'h558; 
        #20 data_in = 12'h559; 
        #20 data_in = 12'h55a; 
        #20 data_in = 12'h55b; 
        #20 data_in = 12'h55c; 
        #20 data_in = 12'h55d; 
        #20 data_in = 12'h55e; 
        #20 data_in = 12'h55f; 
        #20 data_in = 12'h560; 
        #20 data_in = 12'h561; 
        #20 data_in = 12'h562; 
        #20 data_in = 12'h563; 
        #20 data_in = 12'h564; 
        #20 data_in = 12'h565; 
        #20 data_in = 12'h566; 
        #20 data_in = 12'h567; 
        #20 data_in = 12'h568; 
        #20 data_in = 12'h569; 
        #20 data_in = 12'h56a; 
        #20 data_in = 12'h56b; 
        #20 data_in = 12'h56c; 
        #20 data_in = 12'h56d; 
        #20 data_in = 12'h56e; 
        #20 data_in = 12'h56f; 
        #20 data_in = 12'h570; 
        #20 data_in = 12'h571; 
        #20 data_in = 12'h572; 
        #20 data_in = 12'h573; 
        #20 data_in = 12'h574; 
        #20 data_in = 12'h575; 
        #20 data_in = 12'h576; 
        #20 data_in = 12'h577; 
        #20 data_in = 12'h578; 
        #20 data_in = 12'h579; 
        #20 data_in = 12'h57a; 
        #20 data_in = 12'h57b; 
        #20 data_in = 12'h57c; 
        #20 data_in = 12'h57d; 
        #20 data_in = 12'h57e; 
        #20 data_in = 12'h57f; 
        #20 data_in = 12'h580; 
        #20 data_in = 12'h581; 
        #20 data_in = 12'h582; 
        #20 data_in = 12'h583; 
        #20 data_in = 12'h584; 
        #20 data_in = 12'h585; 
        #20 data_in = 12'h586; 
        #20 data_in = 12'h587; 
        #20 data_in = 12'h588; 
        #20 data_in = 12'h589; 
        #20 data_in = 12'h58a; 
        #20 data_in = 12'h58b; 
        #20 data_in = 12'h58c; 
        #20 data_in = 12'h58d; 
        #20 data_in = 12'h58e; 
        #20 data_in = 12'h58f; 
        #20 data_in = 12'h590; 
        #20 data_in = 12'h591; 
        #20 data_in = 12'h592; 
        #20 data_in = 12'h593; 
        #20 data_in = 12'h594; 
        #20 data_in = 12'h595; 
        #20 data_in = 12'h596; 
        #20 data_in = 12'h597; 
        #20 data_in = 12'h598; 
        #20 data_in = 12'h599; 
        #20 data_in = 12'h59a; 
        #20 data_in = 12'h59b; 
        #20 data_in = 12'h59c; 
        #20 data_in = 12'h59d; 
        #20 data_in = 12'h59e; 
        #20 data_in = 12'h59f; 
        #20 data_in = 12'h5a0; 
        #20 data_in = 12'h5a1; 
        #20 data_in = 12'h5a2; 
        #20 data_in = 12'h5a3; 
        #20 data_in = 12'h5a4; 
        #20 data_in = 12'h5a5; 
        #20 data_in = 12'h5a6; 
        #20 data_in = 12'h5a7; 
        #20 data_in = 12'h5a8; 
        #20 data_in = 12'h5a9; 
        #20 data_in = 12'h5aa; 
        #20 data_in = 12'h5ab; 
        #20 data_in = 12'h5ac; 
        #20 data_in = 12'h5ad; 
        #20 data_in = 12'h5ae; 
        #20 data_in = 12'h5af; 
        #20 data_in = 12'h5b0; 
        #20 data_in = 12'h5b1; 
        #20 data_in = 12'h5b2; 
        #20 data_in = 12'h5b3; 
        #20 data_in = 12'h5b4; 
        #20 data_in = 12'h5b5; 
        #20 data_in = 12'h5b6; 
        #20 data_in = 12'h5b7; 
        #20 data_in = 12'h5b8; 
        #20 data_in = 12'h5b9; 
        #20 data_in = 12'h5ba; 
        #20 data_in = 12'h5bb; 
        #20 data_in = 12'h5bc; 
        #20 data_in = 12'h5bd; 
        #20 data_in = 12'h5be; 
        #20 data_in = 12'h5bf; 
        #20 data_in = 12'h5c0; 
        #20 data_in = 12'h5c1; 
        #20 data_in = 12'h5c2; 
        #20 data_in = 12'h5c3; 
        #20 data_in = 12'h5c4; 
        #20 data_in = 12'h5c5; 
        #20 data_in = 12'h5c6; 
        #20 data_in = 12'h5c7; 
        #20 data_in = 12'h5c8; 
        #20 data_in = 12'h5c9; 
        #20 data_in = 12'h5ca; 
        #20 data_in = 12'h5cb; 
        #20 data_in = 12'h5cc; 
        #20 data_in = 12'h5cd; 
        #20 data_in = 12'h5ce; 
        #20 data_in = 12'h5cf; 
        #20 data_in = 12'h5d0; 
        #20 data_in = 12'h5d1; 
        #20 data_in = 12'h5d2; 
        #20 data_in = 12'h5d3; 
        #20 data_in = 12'h5d4; 
        #20 data_in = 12'h5d5; 
        #20 data_in = 12'h5d6; 
        #20 data_in = 12'h5d7; 
        #20 data_in = 12'h5d8; 
        #20 data_in = 12'h5d9; 
        #20 data_in = 12'h5da; 
        #20 data_in = 12'h5db; 
        #20 data_in = 12'h5dc; 
        #20 data_in = 12'h5dd; 
        #20 data_in = 12'h5de; 
        #20 data_in = 12'h5df; 
        #20 data_in = 12'h5e0; 
        #20 data_in = 12'h5e1; 
        #20 data_in = 12'h5e2; 
        #20 data_in = 12'h5e3; 
        #20 data_in = 12'h5e4; 
        #20 data_in = 12'h5e5; 
        #20 data_in = 12'h5e6; 
        #20 data_in = 12'h5e7; 
        #20 data_in = 12'h5e8; 
        #20 data_in = 12'h5e9; 
        #20 data_in = 12'h5ea; 
        #20 data_in = 12'h5eb; 
        #20 data_in = 12'h5ec; 
        #20 data_in = 12'h5ed; 
        #20 data_in = 12'h5ee; 
        #20 data_in = 12'h5ef; 
        #20 data_in = 12'h5f0; 
        #20 data_in = 12'h5f1; 
        #20 data_in = 12'h5f2; 
        #20 data_in = 12'h5f3; 
        #20 data_in = 12'h5f4; 
        #20 data_in = 12'h5f5; 
        #20 data_in = 12'h5f6; 
        #20 data_in = 12'h5f7; 
        #20 data_in = 12'h5f8; 
        #20 data_in = 12'h5f9; 
        #20 data_in = 12'h5fa; 
        #20 data_in = 12'h5fb; 
        #20 data_in = 12'h5fc; 
        #20 data_in = 12'h5fd; 
        #20 data_in = 12'h5fe; 
        #20 data_in = 12'h5ff; 
        #20 data_in = 12'h600; 
        #20 data_in = 12'h601; 
        #20 data_in = 12'h602; 
        #20 data_in = 12'h603; 
        #20 data_in = 12'h604; 
        #20 data_in = 12'h605; 
        #20 data_in = 12'h606; 
        #20 data_in = 12'h607; 
        #20 data_in = 12'h608; 
        #20 data_in = 12'h609; 
        #20 data_in = 12'h60a; 
        #20 data_in = 12'h60b; 
        #20 data_in = 12'h60c; 
        #20 data_in = 12'h60d; 
        #20 data_in = 12'h60e; 
        #20 data_in = 12'h60f; 
        #20 data_in = 12'h610; 
        #20 data_in = 12'h611; 
        #20 data_in = 12'h612; 
        #20 data_in = 12'h613; 
        #20 data_in = 12'h614; 
        #20 data_in = 12'h615; 
        #20 data_in = 12'h616; 
        #20 data_in = 12'h617; 
        #20 data_in = 12'h618; 
        #20 data_in = 12'h619; 
        #20 data_in = 12'h61a; 
        #20 data_in = 12'h61b; 
        #20 data_in = 12'h61c; 
        #20 data_in = 12'h61d; 
        #20 data_in = 12'h61e; 
        #20 data_in = 12'h61f; 
        #20 data_in = 12'h620; 
        #20 data_in = 12'h621; 
        #20 data_in = 12'h622; 
        #20 data_in = 12'h623; 
        #20 data_in = 12'h624; 
        #20 data_in = 12'h625; 
        #20 data_in = 12'h626; 
        #20 data_in = 12'h627; 
        #20 data_in = 12'h628; 
        #20 data_in = 12'h629; 
        #20 data_in = 12'h62a; 
        #20 data_in = 12'h62b; 
        #20 data_in = 12'h62c; 
        #20 data_in = 12'h62d; 
        #20 data_in = 12'h62e; 
        #20 data_in = 12'h62f; 
        #20 data_in = 12'h630; 
        #20 data_in = 12'h631; 
        #20 data_in = 12'h632; 
        #20 data_in = 12'h633; 
        #20 data_in = 12'h634; 
        #20 data_in = 12'h635; 
        #20 data_in = 12'h636; 
        #20 data_in = 12'h637; 
        #20 data_in = 12'h638; 
        #20 data_in = 12'h639; 
        #20 data_in = 12'h63a; 
        #20 data_in = 12'h63b; 
        #20 data_in = 12'h63c; 
        #20 data_in = 12'h63d; 
        #20 data_in = 12'h63e; 
        #20 data_in = 12'h63f; 
        #20 data_in = 12'h640; 
        #20 data_in = 12'h641; 
        #20 data_in = 12'h642; 
        #20 data_in = 12'h643; 
        #20 data_in = 12'h644; 
        #20 data_in = 12'h645; 
        #20 data_in = 12'h646; 
        #20 data_in = 12'h647; 
        #20 data_in = 12'h648; 
        #20 data_in = 12'h649; 
        #20 data_in = 12'h64a; 
        #20 data_in = 12'h64b; 
        #20 data_in = 12'h64c; 
        #20 data_in = 12'h64d; 
        #20 data_in = 12'h64e; 
        #20 data_in = 12'h64f; 
        #20 data_in = 12'h650; 
        #20 data_in = 12'h651; 
        #20 data_in = 12'h652; 
        #20 data_in = 12'h653; 
        #20 data_in = 12'h654; 
        #20 data_in = 12'h655; 
        #20 data_in = 12'h656; 
        #20 data_in = 12'h657; 
        #20 data_in = 12'h658; 
        #20 data_in = 12'h659; 
        #20 data_in = 12'h65a; 
        #20 data_in = 12'h65b; 
        #20 data_in = 12'h65c; 
        #20 data_in = 12'h65d; 
        #20 data_in = 12'h65e; 
        #20 data_in = 12'h65f; 
        #20 data_in = 12'h660; 
        #20 data_in = 12'h661; 
        #20 data_in = 12'h662; 
        #20 data_in = 12'h663; 
        #20 data_in = 12'h664; 
        #20 data_in = 12'h665; 
        #20 data_in = 12'h666; 
        #20 data_in = 12'h667; 
        #20 data_in = 12'h668; 
        #20 data_in = 12'h669; 
        #20 data_in = 12'h66a; 
        #20 data_in = 12'h66b; 
        #20 data_in = 12'h66c; 
        #20 data_in = 12'h66d; 
        #20 data_in = 12'h66e; 
        #20 data_in = 12'h66f; 
        #20 data_in = 12'h670; 
        #20 data_in = 12'h671; 
        #20 data_in = 12'h672; 
        #20 data_in = 12'h673; 
        #20 data_in = 12'h674; 
        #20 data_in = 12'h675; 
        #20 data_in = 12'h676; 
        #20 data_in = 12'h677; 
        #20 data_in = 12'h678; 
        #20 data_in = 12'h679; 
        #20 data_in = 12'h67a; 
        #20 data_in = 12'h67b; 
        #20 data_in = 12'h67c; 
        #20 data_in = 12'h67d; 
        #20 data_in = 12'h67e; 
        #20 data_in = 12'h67f; 
        #20 data_in = 12'h680; 
        #20 data_in = 12'h681; 
        #20 data_in = 12'h682; 
        #20 data_in = 12'h683; 
        #20 data_in = 12'h684; 
        #20 data_in = 12'h685; 
        #20 data_in = 12'h686; 
        #20 data_in = 12'h687; 
        #20 data_in = 12'h688; 
        #20 data_in = 12'h689; 
        #20 data_in = 12'h68a; 
        #20 data_in = 12'h68b; 
        #20 data_in = 12'h68c; 
        #20 data_in = 12'h68d; 
        #20 data_in = 12'h68e; 
        #20 data_in = 12'h68f; 
        #20 data_in = 12'h690; 
        #20 data_in = 12'h691; 
        #20 data_in = 12'h692; 
        #20 data_in = 12'h693; 
        #20 data_in = 12'h694; 
        #20 data_in = 12'h695; 
        #20 data_in = 12'h696; 
        #20 data_in = 12'h697; 
        #20 data_in = 12'h698; 
        #20 data_in = 12'h699; 
        #20 data_in = 12'h69a; 
        #20 data_in = 12'h69b; 
        #20 data_in = 12'h69c; 
        #20 data_in = 12'h69d; 
        #20 data_in = 12'h69e; 
        #20 data_in = 12'h69f; 
        #20 data_in = 12'h6a0; 
        #20 data_in = 12'h6a1; 
        #20 data_in = 12'h6a2; 
        #20 data_in = 12'h6a3; 
        #20 data_in = 12'h6a4; 
        #20 data_in = 12'h6a5; 
        #20 data_in = 12'h6a6; 
        #20 data_in = 12'h6a7; 
        #20 data_in = 12'h6a8; 
        #20 data_in = 12'h6a9; 
        #20 data_in = 12'h6aa; 
        #20 data_in = 12'h6ab; 
        #20 data_in = 12'h6ac; 
        #20 data_in = 12'h6ad; 
        #20 data_in = 12'h6ae; 
        #20 data_in = 12'h6af; 
        #20 data_in = 12'h6b0; 
        #20 data_in = 12'h6b1; 
        #20 data_in = 12'h6b2; 
        #20 data_in = 12'h6b3; 
        #20 data_in = 12'h6b4; 
        #20 data_in = 12'h6b5; 
        #20 data_in = 12'h6b6; 
        #20 data_in = 12'h6b7; 
        #20 data_in = 12'h6b8; 
        #20 data_in = 12'h6b9; 
        #20 data_in = 12'h6ba; 
        #20 data_in = 12'h6bb; 
        #20 data_in = 12'h6bc; 
        #20 data_in = 12'h6bd; 
        #20 data_in = 12'h6be; 
        #20 data_in = 12'h6bf; 
        #20 data_in = 12'h6c0; 
        #20 data_in = 12'h6c1; 
        #20 data_in = 12'h6c2; 
        #20 data_in = 12'h6c3; 
        #20 data_in = 12'h6c4; 
        #20 data_in = 12'h6c5; 
        #20 data_in = 12'h6c6; 
        #20 data_in = 12'h6c7; 
        #20 data_in = 12'h6c8; 
        #20 data_in = 12'h6c9; 
        #20 data_in = 12'h6ca; 
        #20 data_in = 12'h6cb; 
        #20 data_in = 12'h6cc; 
        #20 data_in = 12'h6cd; 
        #20 data_in = 12'h6ce; 
        #20 data_in = 12'h6cf; 
        #20 data_in = 12'h6d0; 
        #20 data_in = 12'h6d1; 
        #20 data_in = 12'h6d2; 
        #20 data_in = 12'h6d3; 
        #20 data_in = 12'h6d4; 
        #20 data_in = 12'h6d5; 
        #20 data_in = 12'h6d6; 
        #20 data_in = 12'h6d7; 
        #20 data_in = 12'h6d8; 
        #20 data_in = 12'h6d9; 
        #20 data_in = 12'h6da; 
        #20 data_in = 12'h6db; 
        #20 data_in = 12'h6dc; 
        #20 data_in = 12'h6dd; 
        #20 data_in = 12'h6de; 
        #20 data_in = 12'h6df; 
        #20 data_in = 12'h6e0; 
        #20 data_in = 12'h6e1; 
        #20 data_in = 12'h6e2; 
        #20 data_in = 12'h6e3; 
        #20 data_in = 12'h6e4; 
        #20 data_in = 12'h6e5; 
        #20 data_in = 12'h6e6; 
        #20 data_in = 12'h6e7; 
        #20 data_in = 12'h6e8; 
        #20 data_in = 12'h6e9; 
        #20 data_in = 12'h6ea; 
        #20 data_in = 12'h6eb; 
        #20 data_in = 12'h6ec; 
        #20 data_in = 12'h6ed; 
        #20 data_in = 12'h6ee; 
        #20 data_in = 12'h6ef; 
        #20 data_in = 12'h6f0; 
        #20 data_in = 12'h6f1; 
        #20 data_in = 12'h6f2; 
        #20 data_in = 12'h6f3; 
        #20 data_in = 12'h6f4; 
        #20 data_in = 12'h6f5; 
        #20 data_in = 12'h6f6; 
        #20 data_in = 12'h6f7; 
        #20 data_in = 12'h6f8; 
        #20 data_in = 12'h6f9; 
        #20 data_in = 12'h6fa; 
        #20 data_in = 12'h6fb; 
        #20 data_in = 12'h6fc; 
        #20 data_in = 12'h6fd; 
        #20 data_in = 12'h6fe; 
        #20 data_in = 12'h6ff; 
        #20 data_in = 12'h700; 
        #20 data_in = 12'h701; 
        #20 data_in = 12'h702; 
        #20 data_in = 12'h703; 
        #20 data_in = 12'h704; 
        #20 data_in = 12'h705; 
        #20 data_in = 12'h706; 
        #20 data_in = 12'h707; 
        #20 data_in = 12'h708; 
        #20 data_in = 12'h709; 
        #20 data_in = 12'h70a; 
        #20 data_in = 12'h70b; 
        #20 data_in = 12'h70c; 
        #20 data_in = 12'h70d; 
        #20 data_in = 12'h70e; 
        #20 data_in = 12'h70f; 
        #20 data_in = 12'h710; 
        #20 data_in = 12'h711; 
        #20 data_in = 12'h712; 
        #20 data_in = 12'h713; 
        #20 data_in = 12'h714; 
        #20 data_in = 12'h715; 
        #20 data_in = 12'h716; 
        #20 data_in = 12'h717; 
        #20 data_in = 12'h718; 
        #20 data_in = 12'h719; 
        #20 data_in = 12'h71a; 
        #20 data_in = 12'h71b; 
        #20 data_in = 12'h71c; 
        #20 data_in = 12'h71d; 
        #20 data_in = 12'h71e; 
        #20 data_in = 12'h71f; 
        #20 data_in = 12'h720; 
        #20 data_in = 12'h721; 
        #20 data_in = 12'h722; 
        #20 data_in = 12'h723; 
        #20 data_in = 12'h724; 
        #20 data_in = 12'h725; 
        #20 data_in = 12'h726; 
        #20 data_in = 12'h727; 
        #20 data_in = 12'h728; 
        #20 data_in = 12'h729; 
        #20 data_in = 12'h72a; 
        #20 data_in = 12'h72b; 
        #20 data_in = 12'h72c; 
        #20 data_in = 12'h72d; 
        #20 data_in = 12'h72e; 
        #20 data_in = 12'h72f; 
        #20 data_in = 12'h730; 
        #20 data_in = 12'h731; 
        #20 data_in = 12'h732; 
        #20 data_in = 12'h733; 
        #20 data_in = 12'h734; 
        #20 data_in = 12'h735; 
        #20 data_in = 12'h736; 
        #20 data_in = 12'h737; 
        #20 data_in = 12'h738; 
        #20 data_in = 12'h739; 
        #20 data_in = 12'h73a; 
        #20 data_in = 12'h73b; 
        #20 data_in = 12'h73c; 
        #20 data_in = 12'h73d; 
        #20 data_in = 12'h73e; 
        #20 data_in = 12'h73f; 
        #20 data_in = 12'h740; 
        #20 data_in = 12'h741; 
        #20 data_in = 12'h742; 
        #20 data_in = 12'h743; 
        #20 data_in = 12'h744; 
        #20 data_in = 12'h745; 
        #20 data_in = 12'h746; 
        #20 data_in = 12'h747; 
        #20 data_in = 12'h748; 
        #20 data_in = 12'h749; 
        #20 data_in = 12'h74a; 
        #20 data_in = 12'h74b; 
        #20 data_in = 12'h74c; 
        #20 data_in = 12'h74d; 
        #20 data_in = 12'h74e; 
        #20 data_in = 12'h74f; 
        #20 data_in = 12'h750; 
        #20 data_in = 12'h751; 
        #20 data_in = 12'h752; 
        #20 data_in = 12'h753; 
        #20 data_in = 12'h754; 
        #20 data_in = 12'h755; 
        #20 data_in = 12'h756; 
        #20 data_in = 12'h757; 
        #20 data_in = 12'h758; 
        #20 data_in = 12'h759; 
        #20 data_in = 12'h75a; 
        #20 data_in = 12'h75b; 
        #20 data_in = 12'h75c; 
        #20 data_in = 12'h75d; 
        #20 data_in = 12'h75e; 
        #20 data_in = 12'h75f; 
        #20 data_in = 12'h760; 
        #20 data_in = 12'h761; 
        #20 data_in = 12'h762; 
        #20 data_in = 12'h763; 
        #20 data_in = 12'h764; 
        #20 data_in = 12'h765; 
        #20 data_in = 12'h766; 
        #20 data_in = 12'h767; 
        #20 data_in = 12'h768; 
        #20 data_in = 12'h769; 
        #20 data_in = 12'h76a; 
        #20 data_in = 12'h76b; 
        #20 data_in = 12'h76c; 
        #20 data_in = 12'h76d; 
        #20 data_in = 12'h76e; 
        #20 data_in = 12'h76f; 
        #20 data_in = 12'h770; 
        #20 data_in = 12'h771; 
        #20 data_in = 12'h772; 
        #20 data_in = 12'h773; 
        #20 data_in = 12'h774; 
        #20 data_in = 12'h775; 
        #20 data_in = 12'h776; 
        #20 data_in = 12'h777; 
        #20 data_in = 12'h778; 
        #20 data_in = 12'h779; 
        #20 data_in = 12'h77a; 
        #20 data_in = 12'h77b; 
        #20 data_in = 12'h77c; 
        #20 data_in = 12'h77d; 
        #20 data_in = 12'h77e; 
        #20 data_in = 12'h77f; 
        #20 data_in = 12'h780; 
        #20 data_in = 12'h781; 
        #20 data_in = 12'h782; 
        #20 data_in = 12'h783; 
        #20 data_in = 12'h784; 
        #20 data_in = 12'h785; 
        #20 data_in = 12'h786; 
        #20 data_in = 12'h787; 
        #20 data_in = 12'h788; 
        #20 data_in = 12'h789; 
        #20 data_in = 12'h78a; 
        #20 data_in = 12'h78b; 
        #20 data_in = 12'h78c; 
        #20 data_in = 12'h78d; 
        #20 data_in = 12'h78e; 
        #20 data_in = 12'h78f; 
        #20 data_in = 12'h790; 
        #20 data_in = 12'h791; 
        #20 data_in = 12'h792; 
        #20 data_in = 12'h793; 
        #20 data_in = 12'h794; 
        #20 data_in = 12'h795; 
        #20 data_in = 12'h796; 
        #20 data_in = 12'h797; 
        #20 data_in = 12'h798; 
        #20 data_in = 12'h799; 
        #20 data_in = 12'h79a; 
        #20 data_in = 12'h79b; 
        #20 data_in = 12'h79c; 
        #20 data_in = 12'h79d; 
        #20 data_in = 12'h79e; 
        #20 data_in = 12'h79f; 
        #20 data_in = 12'h7a0; 
        #20 data_in = 12'h7a1; 
        #20 data_in = 12'h7a2; 
        #20 data_in = 12'h7a3; 
        #20 data_in = 12'h7a4; 
        #20 data_in = 12'h7a5; 
        #20 data_in = 12'h7a6; 
        #20 data_in = 12'h7a7; 
        #20 data_in = 12'h7a8; 
        #20 data_in = 12'h7a9; 
        #20 data_in = 12'h7aa; 
        #20 data_in = 12'h7ab; 
        #20 data_in = 12'h7ac; 
        #20 data_in = 12'h7ad; 
        #20 data_in = 12'h7ae; 
        #20 data_in = 12'h7af; 
        #20 data_in = 12'h7b0; 
        #20 data_in = 12'h7b1; 
        #20 data_in = 12'h7b2; 
        #20 data_in = 12'h7b3; 
        #20 data_in = 12'h7b4; 
        #20 data_in = 12'h7b5; 
        #20 data_in = 12'h7b6; 
        #20 data_in = 12'h7b7; 
        #20 data_in = 12'h7b8; 
        #20 data_in = 12'h7b9; 
        #20 data_in = 12'h7ba; 
        #20 data_in = 12'h7bb; 
        #20 data_in = 12'h7bc; 
        #20 data_in = 12'h7bd; 
        #20 data_in = 12'h7be; 
        #20 data_in = 12'h7bf; 
        #20 data_in = 12'h7c0; 
        #20 data_in = 12'h7c1; 
        #20 data_in = 12'h7c2; 
        #20 data_in = 12'h7c3; 
        #20 data_in = 12'h7c4; 
        #20 data_in = 12'h7c5; 
        #20 data_in = 12'h7c6; 
        #20 data_in = 12'h7c7; 
        #20 data_in = 12'h7c8; 
        #20 data_in = 12'h7c9; 
        #20 data_in = 12'h7ca; 
        #20 data_in = 12'h7cb; 
        #20 data_in = 12'h7cc; 
        #20 data_in = 12'h7cd; 
        #20 data_in = 12'h7ce; 
        #20 data_in = 12'h7cf; 
        #20 data_in = 12'h7d0; 
        #20 data_in = 12'h7d1; 
        #20 data_in = 12'h7d2; 
        #20 data_in = 12'h7d3; 
        #20 data_in = 12'h7d4; 
        #20 data_in = 12'h7d5; 
        #20 data_in = 12'h7d6; 
        #20 data_in = 12'h7d7; 
        #20 data_in = 12'h7d8; 
        #20 data_in = 12'h7d9; 
        #20 data_in = 12'h7da; 
        #20 data_in = 12'h7db; 
        #20 data_in = 12'h7dc; 
        #20 data_in = 12'h7dd; 
        #20 data_in = 12'h7de; 
        #20 data_in = 12'h7df; 
        #20 data_in = 12'h7e0; 
        #20 data_in = 12'h7e1; 
        #20 data_in = 12'h7e2; 
        #20 data_in = 12'h7e3; 
        #20 data_in = 12'h7e4; 
        #20 data_in = 12'h7e5; 
        #20 data_in = 12'h7e6; 
        #20 data_in = 12'h7e7; 
        #20 data_in = 12'h7e8; 
        #20 data_in = 12'h7e9; 
        #20 data_in = 12'h7ea; 
        #20 data_in = 12'h7eb; 
        #20 data_in = 12'h7ec; 
        #20 data_in = 12'h7ed; 
        #20 data_in = 12'h7ee; 
        #20 data_in = 12'h7ef; 
        #20 data_in = 12'h7f0; 
        #20 data_in = 12'h7f1; 
        #20 data_in = 12'h7f2; 
        #20 data_in = 12'h7f3; 
        #20 data_in = 12'h7f4; 
        #20 data_in = 12'h7f5; 
        #20 data_in = 12'h7f6; 
        #20 data_in = 12'h7f7; 
        #20 data_in = 12'h7f8;		
        #20 data_in = 12'h7f9; 
        #20 data_in = 12'h7fa; 
        #20 data_in = 12'h7fb; 
        #20 data_in = 12'h7fc; 
        #20 data_in = 12'h7fd;
        #20 data_in = 12'h7fe; 
        #20 data_in = 12'h7ff;
        #20 data_in = 12'h800;
        #20 data_in = 12'h801; 
        #20 data_in = 12'h802; 
        #20 data_in = 12'h803; 
        #20 data_in = 12'h804; 
        #20 data_in = 12'h805; 
        #20 data_in = 12'h806; 
        #20 data_in = 12'h807; 
        #20 data_in = 12'h808; 
        #20 data_in = 12'h809; 
        #20 data_in = 12'h80a; 
        #20 data_in = 12'h80b; 
        #20 data_in = 12'h80c; 
        #20 data_in = 12'h80d; 
        #20 data_in = 12'h80e; 
        #20 data_in = 12'h80f; 
        #20 data_in = 12'h810; 
        #20 data_in = 12'h811; 
        #20 data_in = 12'h812; 
        #20 data_in = 12'h813; 
        #20 data_in = 12'h814; 
        #20 data_in = 12'h815; 
        #20 data_in = 12'h816; 
        #20 data_in = 12'h817; 
        #20 data_in = 12'h818; 
        #20 data_in = 12'h819; 
        #20 data_in = 12'h81a; 
        #20 data_in = 12'h81b; 
        #20 data_in = 12'h81c; 
        #20 data_in = 12'h81d; 
        #20 data_in = 12'h81e; 
        #20 data_in = 12'h81f; 
        #20 data_in = 12'h820; 
        #20 data_in = 12'h821; 
        #20 data_in = 12'h822; 
        #20 data_in = 12'h823; 
        #20 data_in = 12'h824; 
        #20 data_in = 12'h825; 
        #20 data_in = 12'h826; 
        #20 data_in = 12'h827; 
        #20 data_in = 12'h828; 
        #20 data_in = 12'h829; 
        #20 data_in = 12'h82a; 
        #20 data_in = 12'h82b; 
        #20 data_in = 12'h82c; 
        #20 data_in = 12'h82d; 
        #20 data_in = 12'h82e; 
        #20 data_in = 12'h82f; 
        #20 data_in = 12'h830; 
        #20 data_in = 12'h831; 
        #20 data_in = 12'h832; 
        #20 data_in = 12'h833; 
        #20 data_in = 12'h834; 
        #20 data_in = 12'h835; 
        #20 data_in = 12'h836; 
        #20 data_in = 12'h837; 
        #20 data_in = 12'h838; 
        #20 data_in = 12'h839; 
        #20 data_in = 12'h83a; 
        #20 data_in = 12'h83b; 
        #20 data_in = 12'h83c; 
        #20 data_in = 12'h83d; 
        #20 data_in = 12'h83e; 
        #20 data_in = 12'h83f; 
        #20 data_in = 12'h840; 
        #20 data_in = 12'h841; 
        #20 data_in = 12'h842; 
        #20 data_in = 12'h843; 
        #20 data_in = 12'h844; 
        #20 data_in = 12'h845; 
        #20 data_in = 12'h846; 
        #20 data_in = 12'h847; 
        #20 data_in = 12'h848; 
        #20 data_in = 12'h849; 
        #20 data_in = 12'h84a; 
        #20 data_in = 12'h84b; 
        #20 data_in = 12'h84c; 
        #20 data_in = 12'h84d; 
        #20 data_in = 12'h84e; 
        #20 data_in = 12'h84f; 
        #20 data_in = 12'h850; 
        #20 data_in = 12'h851; 
        #20 data_in = 12'h852; 
        #20 data_in = 12'h853; 
        #20 data_in = 12'h854; 
        #20 data_in = 12'h855; 
        #20 data_in = 12'h856; 
        #20 data_in = 12'h857; 
        #20 data_in = 12'h858; 
        #20 data_in = 12'h859; 
        #20 data_in = 12'h85a; 
        #20 data_in = 12'h85b; 
        #20 data_in = 12'h85c; 
        #20 data_in = 12'h85d; 
        #20 data_in = 12'h85e; 
        #20 data_in = 12'h85f; 
        #20 data_in = 12'h860; 
        #20 data_in = 12'h861; 
        #20 data_in = 12'h862; 
        #20 data_in = 12'h863; 
        #20 data_in = 12'h864; 
        #20 data_in = 12'h865; 
        #20 data_in = 12'h866; 
        #20 data_in = 12'h867; 
        #20 data_in = 12'h868; 
        #20 data_in = 12'h869; 
        #20 data_in = 12'h86a; 
        #20 data_in = 12'h86b; 
        #20 data_in = 12'h86c; 
        #20 data_in = 12'h86d; 
        #20 data_in = 12'h86e; 
        #20 data_in = 12'h86f; 
        #20 data_in = 12'h870; 
        #20 data_in = 12'h871; 
        #20 data_in = 12'h872; 
        #20 data_in = 12'h873; 
        #20 data_in = 12'h874; 
        #20 data_in = 12'h875; 
        #20 data_in = 12'h876; 
        #20 data_in = 12'h877; 
        #20 data_in = 12'h878; 
        #20 data_in = 12'h879; 
        #20 data_in = 12'h87a; 
        #20 data_in = 12'h87b; 
        #20 data_in = 12'h87c; 
        #20 data_in = 12'h87d; 
        #20 data_in = 12'h87e; 
        #20 data_in = 12'h87f; 
        #20 data_in = 12'h880; 
        #20 data_in = 12'h881; 
        #20 data_in = 12'h882; 
        #20 data_in = 12'h883; 
        #20 data_in = 12'h884; 
        #20 data_in = 12'h885; 
        #20 data_in = 12'h886; 
        #20 data_in = 12'h887; 
        #20 data_in = 12'h888; 
        #20 data_in = 12'h889; 
        #20 data_in = 12'h88a; 
        #20 data_in = 12'h88b; 
        #20 data_in = 12'h88c; 
        #20 data_in = 12'h88d; 
        #20 data_in = 12'h88e; 
        #20 data_in = 12'h88f; 
        #20 data_in = 12'h890; 
        #20 data_in = 12'h891; 
        #20 data_in = 12'h892; 
        #20 data_in = 12'h893; 
        #20 data_in = 12'h894; 
        #20 data_in = 12'h895; 
        #20 data_in = 12'h896; 
        #20 data_in = 12'h897; 
        #20 data_in = 12'h898; 
        #20 data_in = 12'h899; 
        #20 data_in = 12'h89a; 
        #20 data_in = 12'h89b; 
        #20 data_in = 12'h89c; 
        #20 data_in = 12'h89d; 
        #20 data_in = 12'h89e; 
        #20 data_in = 12'h89f; 
        #20 data_in = 12'h8a0; 
        #20 data_in = 12'h8a1; 
        #20 data_in = 12'h8a2; 
        #20 data_in = 12'h8a3; 
        #20 data_in = 12'h8a4; 
        #20 data_in = 12'h8a5; 
        #20 data_in = 12'h8a6; 
        #20 data_in = 12'h8a7; 
        #20 data_in = 12'h8a8; 
        #20 data_in = 12'h8a9; 
        #20 data_in = 12'h8aa; 
        #20 data_in = 12'h8ab; 
        #20 data_in = 12'h8ac; 
        #20 data_in = 12'h8ad; 
        #20 data_in = 12'h8ae; 
        #20 data_in = 12'h8af; 
        #20 data_in = 12'h8b0; 
        #20 data_in = 12'h8b1; 
        #20 data_in = 12'h8b2; 
        #20 data_in = 12'h8b3; 
        #20 data_in = 12'h8b4; 
        #20 data_in = 12'h8b5; 
        #20 data_in = 12'h8b6; 
        #20 data_in = 12'h8b7; 
        #20 data_in = 12'h8b8; 
        #20 data_in = 12'h8b9; 
        #20 data_in = 12'h8ba; 
        #20 data_in = 12'h8bb; 
        #20 data_in = 12'h8bc; 
        #20 data_in = 12'h8bd; 
        #20 data_in = 12'h8be; 
        #20 data_in = 12'h8bf; 
        #20 data_in = 12'h8c0; 
        #20 data_in = 12'h8c1; 
        #20 data_in = 12'h8c2; 
        #20 data_in = 12'h8c3; 
        #20 data_in = 12'h8c4; 
        #20 data_in = 12'h8c5; 
        #20 data_in = 12'h8c6; 
        #20 data_in = 12'h8c7; 
        #20 data_in = 12'h8c8; 
        #20 data_in = 12'h8c9; 
        #20 data_in = 12'h8ca; 
        #20 data_in = 12'h8cb; 
        #20 data_in = 12'h8cc; 
        #20 data_in = 12'h8cd; 
        #20 data_in = 12'h8ce; 
        #20 data_in = 12'h8cf; 
        #20 data_in = 12'h8d0; 
        #20 data_in = 12'h8d1; 
        #20 data_in = 12'h8d2; 
        #20 data_in = 12'h8d3; 
        #20 data_in = 12'h8d4; 
        #20 data_in = 12'h8d5; 
        #20 data_in = 12'h8d6; 
        #20 data_in = 12'h8d7; 
        #20 data_in = 12'h8d8; 
        #20 data_in = 12'h8d9; 
        #20 data_in = 12'h8da; 
        #20 data_in = 12'h8db; 
        #20 data_in = 12'h8dc; 
        #20 data_in = 12'h8dd; 
        #20 data_in = 12'h8de; 
        #20 data_in = 12'h8df; 
        #20 data_in = 12'h8e0; 
        #20 data_in = 12'h8e1; 
        #20 data_in = 12'h8e2; 
        #20 data_in = 12'h8e3; 
        #20 data_in = 12'h8e4; 
        #20 data_in = 12'h8e5; 
        #20 data_in = 12'h8e6; 
        #20 data_in = 12'h8e7; 
        #20 data_in = 12'h8e8; 
        #20 data_in = 12'h8e9; 
        #20 data_in = 12'h8ea; 
        #20 data_in = 12'h8eb; 
        #20 data_in = 12'h8ec; 
        #20 data_in = 12'h8ed; 
        #20 data_in = 12'h8ee; 
        #20 data_in = 12'h8ef; 
        #20 data_in = 12'h8f0; 
        #20 data_in = 12'h8f1; 
        #20 data_in = 12'h8f2; 
        #20 data_in = 12'h8f3; 
        #20 data_in = 12'h8f4; 
        #20 data_in = 12'h8f5; 
        #20 data_in = 12'h8f6; 
        #20 data_in = 12'h8f7; 
        #20 data_in = 12'h8f8; 
        #20 data_in = 12'h8f9; 
        #20 data_in = 12'h8fa; 
        #20 data_in = 12'h8fb; 
        #20 data_in = 12'h8fc; 
        #20 data_in = 12'h8fd; 
        #20 data_in = 12'h8fe; 
        #20 data_in = 12'h8ff; 
        #20 data_in = 12'h900; 
        #20 data_in = 12'h901; 
        #20 data_in = 12'h902; 
        #20 data_in = 12'h903; 
        #20 data_in = 12'h904; 
        #20 data_in = 12'h905; 
        #20 data_in = 12'h906; 
        #20 data_in = 12'h907; 
        #20 data_in = 12'h908; 
        #20 data_in = 12'h909; 
        #20 data_in = 12'h90a; 
        #20 data_in = 12'h90b; 
        #20 data_in = 12'h90c; 
        #20 data_in = 12'h90d; 
        #20 data_in = 12'h90e; 
        #20 data_in = 12'h90f; 
        #20 data_in = 12'h910; 
        #20 data_in = 12'h911; 
        #20 data_in = 12'h912; 
        #20 data_in = 12'h913; 
        #20 data_in = 12'h914; 
        #20 data_in = 12'h915; 
        #20 data_in = 12'h916; 
        #20 data_in = 12'h917; 
        #20 data_in = 12'h918; 
        #20 data_in = 12'h919; 
        #20 data_in = 12'h91a; 
        #20 data_in = 12'h91b; 
        #20 data_in = 12'h91c; 
        #20 data_in = 12'h91d; 
        #20 data_in = 12'h91e; 
        #20 data_in = 12'h91f; 
        #20 data_in = 12'h920; 
        #20 data_in = 12'h921; 
        #20 data_in = 12'h922; 
        #20 data_in = 12'h923; 
        #20 data_in = 12'h924; 
        #20 data_in = 12'h925; 
        #20 data_in = 12'h926; 
        #20 data_in = 12'h927; 
        #20 data_in = 12'h928; 
        #20 data_in = 12'h929; 
        #20 data_in = 12'h92a; 
        #20 data_in = 12'h92b; 
        #20 data_in = 12'h92c; 
        #20 data_in = 12'h92d; 
        #20 data_in = 12'h92e; 
        #20 data_in = 12'h92f; 
        #20 data_in = 12'h930; 
        #20 data_in = 12'h931; 
        #20 data_in = 12'h932; 
        #20 data_in = 12'h933; 
        #20 data_in = 12'h934; 
        #20 data_in = 12'h935; 
        #20 data_in = 12'h936; 
        #20 data_in = 12'h937; 
        #20 data_in = 12'h938; 
        #20 data_in = 12'h939; 
        #20 data_in = 12'h93a; 
        #20 data_in = 12'h93b; 
        #20 data_in = 12'h93c; 
        #20 data_in = 12'h93d; 
        #20 data_in = 12'h93e; 
        #20 data_in = 12'h93f; 
        #20 data_in = 12'h940; 
        #20 data_in = 12'h941; 
        #20 data_in = 12'h942; 
        #20 data_in = 12'h943; 
        #20 data_in = 12'h944; 
        #20 data_in = 12'h945; 
        #20 data_in = 12'h946; 
        #20 data_in = 12'h947; 
        #20 data_in = 12'h948; 
        #20 data_in = 12'h949; 
        #20 data_in = 12'h94a; 
        #20 data_in = 12'h94b; 
        #20 data_in = 12'h94c; 
        #20 data_in = 12'h94d; 
        #20 data_in = 12'h94e; 
        #20 data_in = 12'h94f; 
        #20 data_in = 12'h950; 
        #20 data_in = 12'h951; 
        #20 data_in = 12'h952; 
        #20 data_in = 12'h953; 
        #20 data_in = 12'h954; 
        #20 data_in = 12'h955; 
        #20 data_in = 12'h956; 
        #20 data_in = 12'h957; 
        #20 data_in = 12'h958; 
        #20 data_in = 12'h959; 
        #20 data_in = 12'h95a; 
        #20 data_in = 12'h95b; 
        #20 data_in = 12'h95c; 
        #20 data_in = 12'h95d; 
        #20 data_in = 12'h95e; 
        #20 data_in = 12'h95f; 
        #20 data_in = 12'h960; 
        #20 data_in = 12'h961; 
        #20 data_in = 12'h962; 
        #20 data_in = 12'h963; 
        #20 data_in = 12'h964; 
        #20 data_in = 12'h965; 
        #20 data_in = 12'h966; 
        #20 data_in = 12'h967; 
        #20 data_in = 12'h968; 
        #20 data_in = 12'h969; 
        #20 data_in = 12'h96a; 
        #20 data_in = 12'h96b; 
        #20 data_in = 12'h96c; 
        #20 data_in = 12'h96d; 
        #20 data_in = 12'h96e; 
        #20 data_in = 12'h96f; 
        #20 data_in = 12'h970; 
        #20 data_in = 12'h971; 
        #20 data_in = 12'h972; 
        #20 data_in = 12'h973; 
        #20 data_in = 12'h974; 
        #20 data_in = 12'h975; 
        #20 data_in = 12'h976; 
        #20 data_in = 12'h977; 
        #20 data_in = 12'h978; 
        #20 data_in = 12'h979; 
        #20 data_in = 12'h97a; 
        #20 data_in = 12'h97b; 
        #20 data_in = 12'h97c; 
        #20 data_in = 12'h97d; 
        #20 data_in = 12'h97e; 
        #20 data_in = 12'h97f; 
        #20 data_in = 12'h980; 
        #20 data_in = 12'h981; 
        #20 data_in = 12'h982; 
        #20 data_in = 12'h983; 
        #20 data_in = 12'h984; 
        #20 data_in = 12'h985; 
        #20 data_in = 12'h986; 
        #20 data_in = 12'h987; 
        #20 data_in = 12'h988; 
        #20 data_in = 12'h989; 
        #20 data_in = 12'h98a; 
        #20 data_in = 12'h98b; 
        #20 data_in = 12'h98c; 
        #20 data_in = 12'h98d; 
        #20 data_in = 12'h98e; 
        #20 data_in = 12'h98f; 
        #20 data_in = 12'h990; 
        #20 data_in = 12'h991; 
        #20 data_in = 12'h992; 
        #20 data_in = 12'h993; 
        #20 data_in = 12'h994; 
        #20 data_in = 12'h995; 
        #20 data_in = 12'h996; 
        #20 data_in = 12'h997; 
        #20 data_in = 12'h998; 
        #20 data_in = 12'h999; 
        #20 data_in = 12'h99a; 
        #20 data_in = 12'h99b; 
        #20 data_in = 12'h99c; 
        #20 data_in = 12'h99d; 
        #20 data_in = 12'h99e; 
        #20 data_in = 12'h99f; 
        #20 data_in = 12'h9a0; 
        #20 data_in = 12'h9a1; 
        #20 data_in = 12'h9a2; 
        #20 data_in = 12'h9a3; 
        #20 data_in = 12'h9a4; 
        #20 data_in = 12'h9a5; 
        #20 data_in = 12'h9a6; 
        #20 data_in = 12'h9a7; 
        #20 data_in = 12'h9a8; 
        #20 data_in = 12'h9a9; 
        #20 data_in = 12'h9aa; 
        #20 data_in = 12'h9ab; 
        #20 data_in = 12'h9ac; 
        #20 data_in = 12'h9ad; 
        #20 data_in = 12'h9ae; 
        #20 data_in = 12'h9af; 
        #20 data_in = 12'h9b0; 
        #20 data_in = 12'h9b1; 
        #20 data_in = 12'h9b2; 
        #20 data_in = 12'h9b3; 
        #20 data_in = 12'h9b4; 
        #20 data_in = 12'h9b5; 
        #20 data_in = 12'h9b6; 
        #20 data_in = 12'h9b7; 
        #20 data_in = 12'h9b8; 
        #20 data_in = 12'h9b9; 
        #20 data_in = 12'h9ba; 
        #20 data_in = 12'h9bb; 
        #20 data_in = 12'h9bc; 
        #20 data_in = 12'h9bd; 
        #20 data_in = 12'h9be; 
        #20 data_in = 12'h9bf; 
        #20 data_in = 12'h9c0; 
        #20 data_in = 12'h9c1; 
        #20 data_in = 12'h9c2; 
        #20 data_in = 12'h9c3; 
        #20 data_in = 12'h9c4; 
        #20 data_in = 12'h9c5; 
        #20 data_in = 12'h9c6; 
        #20 data_in = 12'h9c7; 
        #20 data_in = 12'h9c8; 
        #20 data_in = 12'h9c9; 
        #20 data_in = 12'h9ca; 
        #20 data_in = 12'h9cb; 
        #20 data_in = 12'h9cc; 
        #20 data_in = 12'h9cd; 
        #20 data_in = 12'h9ce; 
        #20 data_in = 12'h9cf; 
        #20 data_in = 12'h9d0; 
        #20 data_in = 12'h9d1; 
        #20 data_in = 12'h9d2; 
        #20 data_in = 12'h9d3; 
        #20 data_in = 12'h9d4; 
        #20 data_in = 12'h9d5; 
        #20 data_in = 12'h9d6; 
        #20 data_in = 12'h9d7; 
        #20 data_in = 12'h9d8; 
        #20 data_in = 12'h9d9; 
        #20 data_in = 12'h9da; 
        #20 data_in = 12'h9db; 
        #20 data_in = 12'h9dc; 
        #20 data_in = 12'h9dd; 
        #20 data_in = 12'h9de; 
        #20 data_in = 12'h9df; 
        #20 data_in = 12'h9e0; 
        #20 data_in = 12'h9e1; 
        #20 data_in = 12'h9e2; 
        #20 data_in = 12'h9e3; 
        #20 data_in = 12'h9e4; 
        #20 data_in = 12'h9e5; 
        #20 data_in = 12'h9e6; 
        #20 data_in = 12'h9e7; 
        #20 data_in = 12'h9e8; 
        #20 data_in = 12'h9e9; 
        #20 data_in = 12'h9ea; 
        #20 data_in = 12'h9eb; 
        #20 data_in = 12'h9ec; 
        #20 data_in = 12'h9ed; 
        #20 data_in = 12'h9ee; 
        #20 data_in = 12'h9ef; 
        #20 data_in = 12'h9f0; 
        #20 data_in = 12'h9f1; 
        #20 data_in = 12'h9f2; 
        #20 data_in = 12'h9f3; 
        #20 data_in = 12'h9f4; 
        #20 data_in = 12'h9f5; 
        #20 data_in = 12'h9f6; 
        #20 data_in = 12'h9f7; 
        #20 data_in = 12'h9f8; 
        #20 data_in = 12'h9f9; 
        #20 data_in = 12'h9fa; 
        #20 data_in = 12'h9fb; 
        #20 data_in = 12'h9fc; 
        #20 data_in = 12'h9fd; 
        #20 data_in = 12'h9fe; 
        #20 data_in = 12'h9ff; 
        #20 data_in = 12'ha00; 
        #20 data_in = 12'ha01; 
        #20 data_in = 12'ha02; 
        #20 data_in = 12'ha03; 
        #20 data_in = 12'ha04; 
        #20 data_in = 12'ha05; 
        #20 data_in = 12'ha06; 
        #20 data_in = 12'ha07; 
        #20 data_in = 12'ha08; 
        #20 data_in = 12'ha09; 
        #20 data_in = 12'ha0a; 
        #20 data_in = 12'ha0b; 
        #20 data_in = 12'ha0c; 
        #20 data_in = 12'ha0d; 
        #20 data_in = 12'ha0e; 
        #20 data_in = 12'ha0f; 
        #20 data_in = 12'ha10; 
        #20 data_in = 12'ha11; 
        #20 data_in = 12'ha12; 
        #20 data_in = 12'ha13; 
        #20 data_in = 12'ha14; 
        #20 data_in = 12'ha15; 
        #20 data_in = 12'ha16; 
        #20 data_in = 12'ha17; 
        #20 data_in = 12'ha18; 
        #20 data_in = 12'ha19; 
        #20 data_in = 12'ha1a; 
        #20 data_in = 12'ha1b; 
        #20 data_in = 12'ha1c; 
        #20 data_in = 12'ha1d; 
        #20 data_in = 12'ha1e; 
        #20 data_in = 12'ha1f; 
        #20 data_in = 12'ha20; 
        #20 data_in = 12'ha21; 
        #20 data_in = 12'ha22; 
        #20 data_in = 12'ha23; 
        #20 data_in = 12'ha24; 
        #20 data_in = 12'ha25; 
        #20 data_in = 12'ha26; 
        #20 data_in = 12'ha27; 
        #20 data_in = 12'ha28; 
        #20 data_in = 12'ha29; 
        #20 data_in = 12'ha2a; 
        #20 data_in = 12'ha2b; 
        #20 data_in = 12'ha2c; 
        #20 data_in = 12'ha2d; 
        #20 data_in = 12'ha2e; 
        #20 data_in = 12'ha2f; 
        #20 data_in = 12'ha30; 
        #20 data_in = 12'ha31; 
        #20 data_in = 12'ha32; 
        #20 data_in = 12'ha33; 
        #20 data_in = 12'ha34; 
        #20 data_in = 12'ha35; 
        #20 data_in = 12'ha36; 
        #20 data_in = 12'ha37; 
        #20 data_in = 12'ha38; 
        #20 data_in = 12'ha39; 
        #20 data_in = 12'ha3a; 
        #20 data_in = 12'ha3b; 
        #20 data_in = 12'ha3c; 
        #20 data_in = 12'ha3d; 
        #20 data_in = 12'ha3e; 
        #20 data_in = 12'ha3f; 
        #20 data_in = 12'ha40; 
        #20 data_in = 12'ha41; 
        #20 data_in = 12'ha42; 
        #20 data_in = 12'ha43; 
        #20 data_in = 12'ha44; 
        #20 data_in = 12'ha45; 
        #20 data_in = 12'ha46; 
        #20 data_in = 12'ha47; 
        #20 data_in = 12'ha48; 
        #20 data_in = 12'ha49; 
        #20 data_in = 12'ha4a; 
        #20 data_in = 12'ha4b; 
        #20 data_in = 12'ha4c; 
        #20 data_in = 12'ha4d; 
        #20 data_in = 12'ha4e; 
        #20 data_in = 12'ha4f; 
        #20 data_in = 12'ha50; 
        #20 data_in = 12'ha51; 
        #20 data_in = 12'ha52; 
        #20 data_in = 12'ha53; 
        #20 data_in = 12'ha54; 
        #20 data_in = 12'ha55; 
        #20 data_in = 12'ha56; 
        #20 data_in = 12'ha57; 
        #20 data_in = 12'ha58; 
        #20 data_in = 12'ha59; 
        #20 data_in = 12'ha5a; 
        #20 data_in = 12'ha5b; 
        #20 data_in = 12'ha5c; 
        #20 data_in = 12'ha5d; 
        #20 data_in = 12'ha5e; 
        #20 data_in = 12'ha5f; 
        #20 data_in = 12'ha60; 
        #20 data_in = 12'ha61; 
        #20 data_in = 12'ha62; 
        #20 data_in = 12'ha63; 
        #20 data_in = 12'ha64; 
        #20 data_in = 12'ha65; 
        #20 data_in = 12'ha66; 
        #20 data_in = 12'ha67; 
        #20 data_in = 12'ha68; 
        #20 data_in = 12'ha69; 
        #20 data_in = 12'ha6a; 
        #20 data_in = 12'ha6b; 
        #20 data_in = 12'ha6c; 
        #20 data_in = 12'ha6d; 
        #20 data_in = 12'ha6e; 
        #20 data_in = 12'ha6f; 
        #20 data_in = 12'ha70; 
        #20 data_in = 12'ha71; 
        #20 data_in = 12'ha72; 
        #20 data_in = 12'ha73; 
        #20 data_in = 12'ha74; 
        #20 data_in = 12'ha75; 
        #20 data_in = 12'ha76; 
        #20 data_in = 12'ha77; 
        #20 data_in = 12'ha78; 
        #20 data_in = 12'ha79; 
        #20 data_in = 12'ha7a; 
        #20 data_in = 12'ha7b; 
        #20 data_in = 12'ha7c; 
        #20 data_in = 12'ha7d; 
        #20 data_in = 12'ha7e; 
        #20 data_in = 12'ha7f; 
        #20 data_in = 12'ha80; 
        #20 data_in = 12'ha81; 
        #20 data_in = 12'ha82; 
        #20 data_in = 12'ha83; 
        #20 data_in = 12'ha84; 
        #20 data_in = 12'ha85; 
        #20 data_in = 12'ha86; 
        #20 data_in = 12'ha87; 
        #20 data_in = 12'ha88; 
        #20 data_in = 12'ha89; 
        #20 data_in = 12'ha8a; 
        #20 data_in = 12'ha8b; 
        #20 data_in = 12'ha8c; 
        #20 data_in = 12'ha8d; 
        #20 data_in = 12'ha8e; 
        #20 data_in = 12'ha8f; 
        #20 data_in = 12'ha90; 
        #20 data_in = 12'ha91; 
        #20 data_in = 12'ha92; 
        #20 data_in = 12'ha93; 
        #20 data_in = 12'ha94; 
        #20 data_in = 12'ha95; 
        #20 data_in = 12'ha96; 
        #20 data_in = 12'ha97; 
        #20 data_in = 12'ha98; 
        #20 data_in = 12'ha99; 
        #20 data_in = 12'ha9a; 
        #20 data_in = 12'ha9b; 
        #20 data_in = 12'ha9c; 
        #20 data_in = 12'ha9d; 
        #20 data_in = 12'ha9e; 
        #20 data_in = 12'ha9f; 
        #20 data_in = 12'haa0; 
        #20 data_in = 12'haa1; 
        #20 data_in = 12'haa2; 
        #20 data_in = 12'haa3; 
        #20 data_in = 12'haa4; 
        #20 data_in = 12'haa5; 
        #20 data_in = 12'haa6; 
        #20 data_in = 12'haa7; 
        #20 data_in = 12'haa8; 
        #20 data_in = 12'haa9; 
        #20 data_in = 12'haaa; 
        #20 data_in = 12'haab; 
        #20 data_in = 12'haac; 
        #20 data_in = 12'haad; 
        #20 data_in = 12'haae; 
        #20 data_in = 12'haaf; 
        #20 data_in = 12'hab0; 
        #20 data_in = 12'hab1; 
        #20 data_in = 12'hab2; 
        #20 data_in = 12'hab3; 
        #20 data_in = 12'hab4; 
        #20 data_in = 12'hab5; 
        #20 data_in = 12'hab6; 
        #20 data_in = 12'hab7; 
        #20 data_in = 12'hab8; 
        #20 data_in = 12'hab9; 
        #20 data_in = 12'haba; 
        #20 data_in = 12'habb; 
        #20 data_in = 12'habc; 
        #20 data_in = 12'habd; 
        #20 data_in = 12'habe; 
        #20 data_in = 12'habf; 
        #20 data_in = 12'hac0; 
        #20 data_in = 12'hac1; 
        #20 data_in = 12'hac2; 
        #20 data_in = 12'hac3; 
        #20 data_in = 12'hac4; 
        #20 data_in = 12'hac5; 
        #20 data_in = 12'hac6; 
        #20 data_in = 12'hac7; 
        #20 data_in = 12'hac8; 
        #20 data_in = 12'hac9; 
        #20 data_in = 12'haca; 
        #20 data_in = 12'hacb; 
        #20 data_in = 12'hacc; 
        #20 data_in = 12'hacd; 
        #20 data_in = 12'hace; 
        #20 data_in = 12'hacf; 
        #20 data_in = 12'had0; 
        #20 data_in = 12'had1; 
        #20 data_in = 12'had2; 
        #20 data_in = 12'had3; 
        #20 data_in = 12'had4; 
        #20 data_in = 12'had5; 
        #20 data_in = 12'had6; 
        #20 data_in = 12'had7; 
        #20 data_in = 12'had8; 
        #20 data_in = 12'had9; 
        #20 data_in = 12'hada; 
        #20 data_in = 12'hadb; 
        #20 data_in = 12'hadc; 
        #20 data_in = 12'hadd; 
        #20 data_in = 12'hade; 
        #20 data_in = 12'hadf; 
        #20 data_in = 12'hae0; 
        #20 data_in = 12'hae1; 
        #20 data_in = 12'hae2; 
        #20 data_in = 12'hae3; 
        #20 data_in = 12'hae4; 
        #20 data_in = 12'hae5; 
        #20 data_in = 12'hae6; 
        #20 data_in = 12'hae7; 
        #20 data_in = 12'hae8; 
        #20 data_in = 12'hae9; 
        #20 data_in = 12'haea; 
        #20 data_in = 12'haeb; 
        #20 data_in = 12'haec; 
        #20 data_in = 12'haed; 
        #20 data_in = 12'haee; 
        #20 data_in = 12'haef; 
        #20 data_in = 12'haf0; 
        #20 data_in = 12'haf1; 
        #20 data_in = 12'haf2; 
        #20 data_in = 12'haf3; 
        #20 data_in = 12'haf4; 
        #20 data_in = 12'haf5; 
        #20 data_in = 12'haf6; 
        #20 data_in = 12'haf7; 
        #20 data_in = 12'haf8; 
        #20 data_in = 12'haf9; 
        #20 data_in = 12'hafa; 
        #20 data_in = 12'hafb; 
        #20 data_in = 12'hafc; 
        #20 data_in = 12'hafd; 
        #20 data_in = 12'hafe; 
        #20 data_in = 12'haff; 
        #20 data_in = 12'hb00; 
        #20 data_in = 12'hb01; 
        #20 data_in = 12'hb02; 
        #20 data_in = 12'hb03; 
        #20 data_in = 12'hb04; 
        #20 data_in = 12'hb05; 
        #20 data_in = 12'hb06; 
        #20 data_in = 12'hb07; 
        #20 data_in = 12'hb08; 
        #20 data_in = 12'hb09; 
        #20 data_in = 12'hb0a; 
        #20 data_in = 12'hb0b; 
        #20 data_in = 12'hb0c; 
        #20 data_in = 12'hb0d; 
        #20 data_in = 12'hb0e; 
        #20 data_in = 12'hb0f; 
        #20 data_in = 12'hb10; 
        #20 data_in = 12'hb11; 
        #20 data_in = 12'hb12; 
        #20 data_in = 12'hb13; 
        #20 data_in = 12'hb14; 
        #20 data_in = 12'hb15; 
        #20 data_in = 12'hb16; 
        #20 data_in = 12'hb17; 
        #20 data_in = 12'hb18; 
        #20 data_in = 12'hb19; 
        #20 data_in = 12'hb1a; 
        #20 data_in = 12'hb1b; 
        #20 data_in = 12'hb1c; 
        #20 data_in = 12'hb1d; 
        #20 data_in = 12'hb1e; 
        #20 data_in = 12'hb1f; 
        #20 data_in = 12'hb20; 
        #20 data_in = 12'hb21; 
        #20 data_in = 12'hb22; 
        #20 data_in = 12'hb23; 
        #20 data_in = 12'hb24; 
        #20 data_in = 12'hb25; 
        #20 data_in = 12'hb26; 
        #20 data_in = 12'hb27; 
        #20 data_in = 12'hb28; 
        #20 data_in = 12'hb29; 
        #20 data_in = 12'hb2a; 
        #20 data_in = 12'hb2b; 
        #20 data_in = 12'hb2c; 
        #20 data_in = 12'hb2d; 
        #20 data_in = 12'hb2e; 
        #20 data_in = 12'hb2f; 
        #20 data_in = 12'hb30; 
        #20 data_in = 12'hb31; 
        #20 data_in = 12'hb32; 
        #20 data_in = 12'hb33; 
        #20 data_in = 12'hb34; 
        #20 data_in = 12'hb35; 
        #20 data_in = 12'hb36; 
        #20 data_in = 12'hb37; 
        #20 data_in = 12'hb38; 
        #20 data_in = 12'hb39; 
        #20 data_in = 12'hb3a; 
        #20 data_in = 12'hb3b; 
        #20 data_in = 12'hb3c; 
        #20 data_in = 12'hb3d; 
        #20 data_in = 12'hb3e; 
        #20 data_in = 12'hb3f; 
        #20 data_in = 12'hb40; 
        #20 data_in = 12'hb41; 
        #20 data_in = 12'hb42; 
        #20 data_in = 12'hb43; 
        #20 data_in = 12'hb44; 
        #20 data_in = 12'hb45; 
        #20 data_in = 12'hb46; 
        #20 data_in = 12'hb47; 
        #20 data_in = 12'hb48; 
        #20 data_in = 12'hb49; 
        #20 data_in = 12'hb4a; 
        #20 data_in = 12'hb4b; 
        #20 data_in = 12'hb4c; 
        #20 data_in = 12'hb4d; 
        #20 data_in = 12'hb4e; 
        #20 data_in = 12'hb4f; 
        #20 data_in = 12'hb50; 
        #20 data_in = 12'hb51; 
        #20 data_in = 12'hb52; 
        #20 data_in = 12'hb53; 
        #20 data_in = 12'hb54; 
        #20 data_in = 12'hb55; 
        #20 data_in = 12'hb56; 
        #20 data_in = 12'hb57; 
        #20 data_in = 12'hb58; 
        #20 data_in = 12'hb59; 
        #20 data_in = 12'hb5a; 
        #20 data_in = 12'hb5b; 
        #20 data_in = 12'hb5c; 
        #20 data_in = 12'hb5d; 
        #20 data_in = 12'hb5e; 
        #20 data_in = 12'hb5f; 
        #20 data_in = 12'hb60; 
        #20 data_in = 12'hb61; 
        #20 data_in = 12'hb62; 
        #20 data_in = 12'hb63; 
        #20 data_in = 12'hb64; 
        #20 data_in = 12'hb65; 
        #20 data_in = 12'hb66; 
        #20 data_in = 12'hb67; 
        #20 data_in = 12'hb68; 
        #20 data_in = 12'hb69; 
        #20 data_in = 12'hb6a; 
        #20 data_in = 12'hb6b; 
        #20 data_in = 12'hb6c; 
        #20 data_in = 12'hb6d; 
        #20 data_in = 12'hb6e; 
        #20 data_in = 12'hb6f; 
        #20 data_in = 12'hb70; 
        #20 data_in = 12'hb71; 
        #20 data_in = 12'hb72; 
        #20 data_in = 12'hb73; 
        #20 data_in = 12'hb74; 
        #20 data_in = 12'hb75; 
        #20 data_in = 12'hb76; 
        #20 data_in = 12'hb77; 
        #20 data_in = 12'hb78; 
        #20 data_in = 12'hb79; 
        #20 data_in = 12'hb7a; 
        #20 data_in = 12'hb7b; 
        #20 data_in = 12'hb7c; 
        #20 data_in = 12'hb7d; 
        #20 data_in = 12'hb7e; 
        #20 data_in = 12'hb7f; 
        #20 data_in = 12'hb80; 
        #20 data_in = 12'hb81; 
        #20 data_in = 12'hb82; 
        #20 data_in = 12'hb83; 
        #20 data_in = 12'hb84; 
        #20 data_in = 12'hb85; 
        #20 data_in = 12'hb86; 
        #20 data_in = 12'hb87; 
        #20 data_in = 12'hb88; 
        #20 data_in = 12'hb89; 
        #20 data_in = 12'hb8a; 
        #20 data_in = 12'hb8b; 
        #20 data_in = 12'hb8c; 
        #20 data_in = 12'hb8d; 
        #20 data_in = 12'hb8e; 
        #20 data_in = 12'hb8f; 
        #20 data_in = 12'hb90; 
        #20 data_in = 12'hb91; 
        #20 data_in = 12'hb92; 
        #20 data_in = 12'hb93; 
        #20 data_in = 12'hb94; 
        #20 data_in = 12'hb95; 
        #20 data_in = 12'hb96; 
        #20 data_in = 12'hb97; 
        #20 data_in = 12'hb98; 
        #20 data_in = 12'hb99; 
        #20 data_in = 12'hb9a; 
        #20 data_in = 12'hb9b; 
        #20 data_in = 12'hb9c; 
        #20 data_in = 12'hb9d; 
        #20 data_in = 12'hb9e; 
        #20 data_in = 12'hb9f; 
        #20 data_in = 12'hba0;	read    = 1;		
        #20 data_in = 12'hba1; 
        #20 data_in = 12'hba2; 
        #20 data_in = 12'hba3; 
        #20 data_in = 12'hba4; 
        #20 data_in = 12'hba5; 
        #20 data_in = 12'hba6; 
        #20 data_in = 12'hba7; 
        #20 data_in = 12'hba8; 
        #20 data_in = 12'hba9; 
        #20 data_in = 12'hbaa;	read    = 0;		
        #20 data_in = 12'hbab; 
        #20 data_in = 12'hbac; 
        #20 data_in = 12'hbad; 
        #20 data_in = 12'hbae; 
        #20 data_in = 12'hbaf; 
        #20 data_in = 12'hbb0;	read    = 1;		
        #20 data_in = 12'hbb1; 
        #20 data_in = 12'hbb2; 
        #20 data_in = 12'hbb3; 
        #20 data_in = 12'hbb4; 
        #20 data_in = 12'hbb5; 
        #20 data_in = 12'hbb6; 
        #20 data_in = 12'hbb7; 
        #20 data_in = 12'hbb8; 	write   = 0;
		#20 $stop;	
    end
endmodule